module top(n0, n1, n2, n3, n4, n5, n6, n7);
    input n0, n1, n2, n3;
    input [15:0] n4;
    output [15:0] n5;
    output n6, n7;
    wire n0, n1, n2, n3;
    wire [15:0] n4;
    wire [15:0] n5;
    wire n6, n7;
    wire [15:0] n8;
    wire [15:0] n9;
    wire [15:0] n10;
    wire [15:0] n11;
    wire [15:0] n12;
    wire [15:0] n13;
    wire [15:0] n14;
    wire [15:0] n15;
    wire [15:0] n16;
    wire [15:0] n17;
    wire [15:0] n18;
    wire [15:0] n19;
    wire [15:0] n20;
    wire [15:0] n21;
    wire [15:0] n22;
    wire [15:0] n23;
    wire [15:0] n24;
    wire [15:0] n25;
    wire [15:0] n26;
    wire [15:0] n27;
    wire [15:0] n28;
    wire [15:0] n29;
    wire [15:0] n30;
    wire n31, n32, n33, n34, n35, n36, n37, n38;
    wire n39, n40, n41, n42, n43, n44, n45, n46;
    wire n47, n48, n49, n50, n51, n52, n53, n54;
    wire n55, n56, n57, n58, n59, n60, n61, n62;
    wire n63, n64, n65, n66, n67, n68, n69, n70;
    wire n71, n72, n73, n74, n75, n76, n77, n78;
    wire n79, n80, n81, n82, n83, n84, n85, n86;
    wire n87, n88, n89, n90, n91, n92, n93, n94;
    wire n95, n96, n97, n98, n99, n100, n101, n102;
    wire n103, n104, n105, n106, n107, n108, n109, n110;
    wire n111, n112, n113, n114, n115, n116, n117, n118;
    wire n119, n120, n121, n122, n123, n124, n125, n126;
    wire n127, n128, n129, n130, n131, n132, n133, n134;
    wire n135, n136, n137, n138, n139, n140, n141, n142;
    wire n143, n144, n145, n146, n147, n148, n149, n150;
    wire n151, n152, n153, n154, n155, n156, n157, n158;
    wire n159, n160, n161, n162, n163, n164, n165, n166;
    wire n167, n168, n169, n170, n171, n172, n173, n174;
    wire n175, n176, n177, n178, n179, n180, n181, n182;
    wire n183, n184, n185, n186, n187, n188, n189, n190;
    wire n191, n192, n193, n194, n195, n196, n197, n198;
    wire n199, n200, n201, n202, n203, n204, n205, n206;
    wire n207, n208, n209, n210, n211, n212, n213, n214;
    wire n215, n216, n217, n218, n219, n220, n221, n222;
    wire n223, n224, n225, n226, n227, n228, n229, n230;
    wire n231, n232, n233, n234, n235, n236, n237, n238;
    wire n239, n240, n241, n242, n243, n244, n245, n246;
    wire n247, n248, n249, n250, n251, n252, n253, n254;
    wire n255, n256, n257, n258, n259, n260, n261, n262;
    wire n263, n264, n265, n266, n267, n268, n269, n270;
    wire n271, n272, n273, n274, n275, n276, n277, n278;
    wire n279, n280, n281, n282, n283, n284, n285, n286;
    wire n287, n288, n289, n290, n291, n292, n293, n294;
    wire n295, n296, n297, n298, n299, n300, n301, n302;
    wire n303, n304, n305, n306, n307, n308, n309, n310;
    wire n311, n312, n313, n314, n315, n316, n317, n318;
    wire n319, n320, n321, n322, n323, n324, n325, n326;
    wire n327, n328, n329, n330, n331, n332, n333, n334;
    wire n335, n336, n337, n338, n339, n340, n341, n342;
    wire n343, n344, n345, n346, n347, n348, n349, n350;
    wire n351, n352, n353, n354, n355, n356, n357, n358;
    wire n359, n360, n361, n362, n363, n364, n365, n366;
    wire n367, n368, n369, n370, n371, n372, n373, n374;
    wire n375, n376, n377, n378, n379, n380, n381, n382;
    wire n383, n384, n385, n386, n387, n388, n389, n390;
    wire n391, n392, n393, n394, n395, n396, n397, n398;
    wire n399, n400, n401, n402, n403, n404, n405, n406;
    wire n407, n408, n409, n410, n411, n412, n413, n414;
    wire n415, n416, n417, n418, n419, n420, n421, n422;
    wire n423, n424, n425, n426, n427, n428, n429, n430;
    wire n431, n432, n433, n434, n435, n436, n437, n438;
    wire n439, n440, n441, n442, n443, n444, n445, n446;
    wire n447, n448, n449, n450, n451, n452, n453, n454;
    wire n455, n456, n457, n458, n459, n460, n461, n462;
    wire n463, n464, n465, n466, n467, n468, n469, n470;
    wire n471, n472, n473, n474, n475, n476, n477, n478;
    wire n479, n480, n481, n482, n483, n484, n485, n486;
    wire n487, n488, n489, n490, n491, n492, n493, n494;
    wire n495, n496, n497, n498, n499, n500, n501, n502;
    wire n503, n504, n505, n506, n507, n508, n509, n510;
    wire n511, n512, n513, n514, n515, n516, n517, n518;
    wire n519, n520, n521, n522, n523, n524, n525, n526;
    wire n527, n528, n529, n530, n531, n532, n533, n534;
    wire n535, n536, n537, n538, n539, n540, n541, n542;
    wire n543, n544, n545, n546, n547, n548, n549, n550;
    wire n551, n552, n553, n554, n555, n556, n557, n558;
    wire n559, n560, n561, n562, n563, n564, n565, n566;
    wire n567, n568, n569, n570, n571, n572, n573, n574;
    wire n575, n576, n577, n578, n579, n580, n581, n582;
    wire n583, n584, n585, n586, n587, n588, n589, n590;
    wire n591, n592, n593, n594, n595, n596, n597, n598;
    wire n599, n600, n601, n602, n603, n604, n605, n606;
    wire n607, n608, n609, n610, n611, n612, n613, n614;
    wire n615, n616, n617, n618, n619, n620, n621, n622;
    wire n623, n624, n625, n626, n627, n628, n629, n630;
    wire n631, n632, n633, n634, n635, n636, n637, n638;
    wire n639, n640, n641, n642, n643, n644, n645, n646;
    wire n647, n648, n649, n650, n651, n652, n653, n654;
    wire n655, n656, n657, n658, n659, n660, n661, n662;
    wire n663, n664, n665, n666, n667, n668, n669, n670;
    wire n671, n672, n673, n674, n675, n676, n677, n678;
    wire n679, n680, n681, n682, n683, n684, n685, n686;
    wire n687, n688, n689, n690, n691, n692, n693, n694;
    wire n695, n696, n697, n698, n699, n700, n701, n702;
    wire n703, n704, n705, n706, n707, n708, n709, n710;
    wire n711, n712, n713, n714, n715, n716, n717, n718;
    wire n719, n720, n721, n722, n723, n724, n725, n726;
    wire n727, n728, n729, n730, n731, n732, n733, n734;
    wire n735, n736, n737, n738, n739, n740, n741, n742;
    wire n743, n744, n745, n746, n747, n748, n749, n750;
    wire n751, n752, n753, n754, n755, n756, n757, n758;
    wire n759, n760, n761, n762, n763, n764, n765, n766;
    wire n767, n768, n769, n770, n771, n772, n773, n774;
    wire n775, n776, n777, n778, n779, n780, n781, n782;
    wire n783, n784, n785, n786, n787, n788, n789, n790;
    wire n791, n792, n793, n794, n795, n796, n797, n798;
    wire n799, n800, n801, n802, n803, n804, n805, n806;
    wire n807, n808, n809, n810, n811, n812, n813, n814;
    wire n815, n816, n817, n818, n819, n820, n821, n822;
    wire n823, n824, n825, n826, n827, n828, n829, n830;
    wire n831, n832, n833, n834, n835, n836, n837, n838;
    wire n839, n840, n841, n842, n843, n844, n845, n846;
    wire n847, n848, n849, n850, n851, n852, n853, n854;
    wire n855, n856, n857, n858, n859, n860, n861, n862;
    wire n863, n864, n865, n866, n867, n868, n869, n870;
    wire n871, n872, n873, n874, n875, n876, n877, n878;
    wire n879, n880, n881, n882, n883, n884, n885, n886;
    wire n887, n888, n889, n890, n891, n892, n893, n894;
    wire n895, n896, n897, n898, n899, n900, n901, n902;
    wire n903, n904, n905, n906, n907, n908, n909, n910;
    wire n911, n912, n913, n914, n915, n916, n917, n918;
    wire n919, n920, n921, n922, n923, n924, n925, n926;
    wire n927, n928, n929, n930, n931, n932, n933, n934;
    wire n935, n936, n937, n938, n939, n940, n941, n942;
    wire n943, n944, n945, n946, n947, n948, n949, n950;
    wire n951, n952, n953, n954, n955, n956, n957, n958;
    wire n959, n960, n961, n962, n963, n964, n965, n966;
    wire n967, n968, n969, n970, n971, n972, n973, n974;
    wire n975, n976, n977, n978, n979, n980, n981, n982;
    wire n983, n984, n985, n986, n987, n988, n989, n990;
    wire n991, n992, n993, n994, n995, n996, n997, n998;
    wire n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006;
    wire n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014;
    wire n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022;
    wire n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030;
    wire n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038;
    wire n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046;
    wire n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054;
    wire n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062;
    wire n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070;
    wire n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078;
    wire n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086;
    wire n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094;
    wire n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102;
    wire n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110;
    wire n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118;
    wire n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126;
    wire n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134;
    wire n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142;
    wire n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150;
    wire n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158;
    wire n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166;
    wire n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174;
    wire n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182;
    wire n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190;
    wire n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198;
    wire n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206;
    wire n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214;
    wire n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222;
    wire n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230;
    wire n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238;
    wire n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246;
    wire n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254;
    wire n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262;
    wire n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270;
    wire n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278;
    wire n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286;
    wire n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294;
    wire n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302;
    wire n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310;
    wire n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318;
    wire n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326;
    wire n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334;
    wire n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342;
    wire n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350;
    wire n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358;
    wire n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366;
    wire n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374;
    wire n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382;
    wire n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390;
    wire n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398;
    wire n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406;
    wire n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414;
    wire n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422;
    wire n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430;
    wire n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438;
    wire n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446;
    wire n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454;
    wire n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462;
    wire n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470;
    wire n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478;
    wire n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486;
    wire n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494;
    wire n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502;
    wire n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510;
    wire n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518;
    wire n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526;
    wire n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534;
    wire n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542;
    wire n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550;
    wire n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558;
    wire n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566;
    wire n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574;
    wire n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582;
    wire n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590;
    wire n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598;
    wire n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606;
    wire n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614;
    wire n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622;
    wire n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630;
    wire n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638;
    wire n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646;
    wire n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654;
    wire n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662;
    wire n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670;
    wire n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678;
    wire n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686;
    wire n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694;
    wire n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702;
    wire n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710;
    wire n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718;
    wire n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726;
    wire n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734;
    wire n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742;
    wire n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750;
    wire n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758;
    wire n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766;
    wire n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774;
    wire n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782;
    wire n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790;
    wire n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798;
    wire n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806;
    wire n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814;
    wire n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822;
    wire n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830;
    wire n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838;
    wire n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846;
    wire n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854;
    wire n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862;
    wire n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870;
    wire n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878;
    wire n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886;
    wire n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894;
    wire n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902;
    wire n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910;
    wire n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918;
    wire n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926;
    wire n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934;
    wire n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942;
    wire n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950;
    wire n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958;
    wire n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966;
    wire n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974;
    wire n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982;
    wire n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990;
    wire n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998;
    wire n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006;
    wire n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014;
    wire n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022;
    wire n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030;
    wire n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038;
    wire n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046;
    wire n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054;
    wire n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062;
    wire n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070;
    wire n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078;
    wire n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086;
    wire n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094;
    wire n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102;
    wire n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110;
    wire n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118;
    wire n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126;
    wire n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134;
    wire n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142;
    wire n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150;
    wire n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158;
    wire n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166;
    wire n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174;
    wire n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182;
    wire n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190;
    wire n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198;
    wire n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206;
    wire n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214;
    wire n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222;
    wire n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230;
    wire n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238;
    wire n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246;
    wire n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254;
    wire n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262;
    wire n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270;
    wire n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278;
    wire n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286;
    wire n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294;
    wire n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302;
    wire n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310;
    wire n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318;
    wire n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326;
    wire n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334;
    wire n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342;
    wire n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350;
    wire n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358;
    wire n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366;
    wire n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374;
    wire n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382;
    wire n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390;
    wire n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398;
    wire n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406;
    wire n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414;
    wire n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422;
    wire n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430;
    wire n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438;
    wire n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446;
    wire n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454;
    wire n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462;
    wire n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470;
    wire n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478;
    wire n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486;
    wire n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494;
    wire n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502;
    wire n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510;
    wire n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518;
    wire n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526;
    wire n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534;
    wire n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542;
    wire n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550;
    wire n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558;
    wire n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566;
    wire n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574;
    wire n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582;
    wire n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590;
    wire n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598;
    wire n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606;
    wire n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614;
    wire n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622;
    wire n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630;
    wire n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638;
    wire n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646;
    wire n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654;
    wire n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662;
    wire n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670;
    wire n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678;
    wire n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686;
    wire n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694;
    wire n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702;
    wire n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710;
    wire n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718;
    wire n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726;
    wire n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734;
    wire n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742;
    wire n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750;
    wire n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758;
    wire n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766;
    wire n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774;
    wire n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782;
    wire n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790;
    wire n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798;
    wire n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806;
    wire n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814;
    wire n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822;
    wire n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830;
    wire n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838;
    wire n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846;
    wire n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854;
    wire n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862;
    wire n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870;
    wire n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878;
    wire n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886;
    wire n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894;
    wire n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902;
    wire n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910;
    wire n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918;
    wire n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926;
    wire n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934;
    wire n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942;
    wire n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950;
    wire n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958;
    wire n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966;
    wire n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974;
    wire n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982;
    wire n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990;
    wire n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998;
    wire n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006;
    wire n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014;
    wire n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022;
    wire n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030;
    wire n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038;
    wire n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046;
    wire n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054;
    wire n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062;
    wire n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070;
    wire n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078;
    wire n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086;
    wire n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094;
    wire n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102;
    wire n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110;
    wire n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118;
    wire n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126;
    wire n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134;
    wire n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142;
    wire n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150;
    wire n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158;
    wire n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166;
    wire n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174;
    wire n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182;
    wire n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190;
    wire n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198;
    wire n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206;
    wire n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214;
    wire n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222;
    wire n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230;
    wire n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238;
    wire n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246;
    wire n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254;
    wire n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262;
    wire n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270;
    wire n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278;
    wire n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286;
    wire n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294;
    wire n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302;
    wire n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310;
    wire n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318;
    wire n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326;
    wire n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334;
    wire n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342;
    wire n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350;
    wire n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358;
    wire n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366;
    wire n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374;
    wire n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382;
    wire n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390;
    wire n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398;
    wire n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406;
    wire n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414;
    wire n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422;
    wire n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430;
    wire n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438;
    wire n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446;
    wire n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454;
    wire n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462;
    wire n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470;
    wire n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478;
    wire n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486;
    wire n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494;
    wire n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502;
    wire n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510;
    wire n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518;
    wire n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526;
    wire n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534;
    wire n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542;
    wire n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550;
    wire n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558;
    wire n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566;
    wire n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574;
    wire n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582;
    wire n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590;
    wire n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598;
    wire n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606;
    wire n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614;
    wire n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622;
    wire n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630;
    wire n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638;
    wire n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646;
    wire n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654;
    wire n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662;
    wire n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670;
    wire n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678;
    wire n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686;
    wire n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694;
    dff g0(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2016), .Q(n6));
    dff g1(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2009), .Q(n7));
    dff g2(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1021), .Q(n24[0]));
    dff g3(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1020), .Q(n24[1]));
    dff g4(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1019), .Q(n24[2]));
    dff g5(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1018), .Q(n24[3]));
    dff g6(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1030), .Q(n25[0]));
    dff g7(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1016), .Q(n25[1]));
    dff g8(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1015), .Q(n25[2]));
    dff g9(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1013), .Q(n25[3]));
    dff g10(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1722), .Q(n26[0]));
    dff g11(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1971), .Q(n26[1]));
    dff g12(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1970), .Q(n26[2]));
    dff g13(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1969), .Q(n26[3]));
    dff g14(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1968), .Q(n26[4]));
    dff g15(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1967), .Q(n26[5]));
    dff g16(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1966), .Q(n26[6]));
    dff g17(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1965), .Q(n26[7]));
    dff g18(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1964), .Q(n26[8]));
    dff g19(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1963), .Q(n26[9]));
    dff g20(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1962), .Q(n26[10]));
    dff g21(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1961), .Q(n26[11]));
    dff g22(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1960), .Q(n26[12]));
    dff g23(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1959), .Q(n26[13]));
    dff g24(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1958), .Q(n26[14]));
    dff g25(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1989), .Q(n26[15]));
    dff g26(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2169), .Q(n5[0]));
    dff g27(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2179), .Q(n5[1]));
    dff g28(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2168), .Q(n5[2]));
    dff g29(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2171), .Q(n5[3]));
    dff g30(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2170), .Q(n5[4]));
    dff g31(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2172), .Q(n5[5]));
    dff g32(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2167), .Q(n5[6]));
    dff g33(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2166), .Q(n5[7]));
    dff g34(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2165), .Q(n5[8]));
    dff g35(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2173), .Q(n5[9]));
    dff g36(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2178), .Q(n5[10]));
    dff g37(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2177), .Q(n5[11]));
    dff g38(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2176), .Q(n5[12]));
    dff g39(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2175), .Q(n5[13]));
    dff g40(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2174), .Q(n5[14]));
    dff g41(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2119), .Q(n5[15]));
    dff g42(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n519), .Q(n27[0]));
    dff g43(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n520), .Q(n27[1]));
    dff g44(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n523), .Q(n27[2]));
    dff g45(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n521), .Q(n27[3]));
    dff g46(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n525), .Q(n28[0]));
    dff g47(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n522), .Q(n28[1]));
    dff g48(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n524), .Q(n28[2]));
    dff g49(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n518), .Q(n28[3]));
    or g50(n2179 ,n2081 ,n2156);
    or g51(n2178 ,n2087 ,n2162);
    or g52(n2177 ,n2086 ,n2161);
    or g53(n2176 ,n2085 ,n2160);
    or g54(n2175 ,n2084 ,n2159);
    or g55(n2174 ,n2083 ,n2164);
    or g56(n2173 ,n2088 ,n2158);
    or g57(n2172 ,n2077 ,n2152);
    or g58(n2171 ,n2079 ,n2154);
    or g59(n2170 ,n2078 ,n2157);
    or g60(n2169 ,n2082 ,n2153);
    or g61(n2168 ,n2080 ,n2155);
    or g62(n2167 ,n2076 ,n2151);
    or g63(n2166 ,n2075 ,n2150);
    or g64(n2165 ,n2074 ,n2163);
    or g65(n2164 ,n627 ,n2145);
    or g66(n2163 ,n630 ,n2148);
    or g67(n2162 ,n633 ,n2146);
    or g68(n2161 ,n625 ,n2149);
    or g69(n2160 ,n624 ,n2144);
    or g70(n2159 ,n632 ,n2143);
    or g71(n2158 ,n631 ,n2147);
    or g72(n2157 ,n621 ,n2142);
    or g73(n2156 ,n622 ,n2141);
    or g74(n2155 ,n623 ,n2140);
    or g75(n2154 ,n636 ,n2139);
    or g76(n2153 ,n626 ,n2138);
    or g77(n2152 ,n635 ,n2137);
    or g78(n2151 ,n628 ,n2136);
    or g79(n2150 ,n629 ,n2135);
    nor g80(n2149 ,n2115 ,n2131);
    nor g81(n2148 ,n2096 ,n2130);
    nor g82(n2147 ,n2117 ,n2133);
    nor g83(n2146 ,n2116 ,n2132);
    nor g84(n2145 ,n2112 ,n2128);
    nor g85(n2144 ,n2114 ,n2134);
    nor g86(n2143 ,n2113 ,n2129);
    nor g87(n2142 ,n2111 ,n2123);
    nor g88(n2141 ,n2106 ,n2122);
    nor g89(n2140 ,n2105 ,n2125);
    nor g90(n2139 ,n2104 ,n2124);
    nor g91(n2138 ,n2107 ,n2127);
    nor g92(n2137 ,n2110 ,n2126);
    nor g93(n2136 ,n2109 ,n2121);
    nor g94(n2135 ,n2108 ,n2120);
    or g95(n2134 ,n785 ,n2099);
    or g96(n2133 ,n785 ,n2102);
    or g97(n2132 ,n785 ,n2101);
    or g98(n2131 ,n785 ,n2100);
    or g99(n2130 ,n785 ,n2103);
    or g100(n2129 ,n785 ,n2098);
    or g101(n2128 ,n785 ,n2097);
    or g102(n2127 ,n785 ,n2118);
    or g103(n2126 ,n785 ,n2091);
    or g104(n2125 ,n785 ,n2094);
    or g105(n2124 ,n785 ,n2093);
    or g106(n2123 ,n785 ,n2092);
    or g107(n2122 ,n785 ,n2073);
    or g108(n2121 ,n785 ,n2090);
    or g109(n2120 ,n785 ,n2089);
    or g110(n2119 ,n634 ,n2095);
    nor g111(n2118 ,n29[0] ,n2060);
    nor g112(n2117 ,n153 ,n2065);
    nor g113(n2116 ,n151 ,n2071);
    nor g114(n2115 ,n147 ,n2069);
    nor g115(n2114 ,n146 ,n2067);
    nor g116(n2113 ,n156 ,n2061);
    nor g117(n2112 ,n150 ,n2063);
    nor g118(n2111 ,n148 ,n2050);
    nor g119(n2110 ,n149 ,n2056);
    nor g120(n2109 ,n155 ,n2046);
    nor g121(n2108 ,n154 ,n2044);
    nor g122(n2107 ,n136 ,n2059);
    nor g123(n2106 ,n139 ,n2048);
    nor g124(n2105 ,n138 ,n2054);
    nor g125(n2104 ,n137 ,n2052);
    nor g126(n2103 ,n29[8] ,n2043);
    nor g127(n2102 ,n29[9] ,n2066);
    nor g128(n2101 ,n29[10] ,n2072);
    nor g129(n2100 ,n29[11] ,n2070);
    nor g130(n2099 ,n29[12] ,n2068);
    nor g131(n2098 ,n29[13] ,n2062);
    nor g132(n2097 ,n29[14] ,n2064);
    nor g133(n2096 ,n145 ,n2042);
    nor g134(n2095 ,n1061 ,n2058);
    nor g135(n2094 ,n29[2] ,n2055);
    nor g136(n2093 ,n29[3] ,n2053);
    nor g137(n2092 ,n29[4] ,n2051);
    nor g138(n2091 ,n29[5] ,n2057);
    nor g139(n2090 ,n29[6] ,n2047);
    nor g140(n2089 ,n29[7] ,n2045);
    nor g141(n2088 ,n783 ,n2065);
    nor g142(n2087 ,n783 ,n2071);
    nor g143(n2086 ,n783 ,n2069);
    nor g144(n2085 ,n783 ,n2067);
    nor g145(n2084 ,n783 ,n2061);
    nor g146(n2083 ,n783 ,n2063);
    nor g147(n2082 ,n783 ,n2059);
    nor g148(n2081 ,n783 ,n2048);
    nor g149(n2080 ,n783 ,n2054);
    nor g150(n2079 ,n783 ,n2052);
    nor g151(n2078 ,n783 ,n2050);
    nor g152(n2077 ,n783 ,n2056);
    nor g153(n2076 ,n783 ,n2046);
    nor g154(n2075 ,n783 ,n2044);
    nor g155(n2074 ,n783 ,n2042);
    nor g156(n2073 ,n29[1] ,n2049);
    not g157(n2072 ,n2071);
    not g158(n2070 ,n2069);
    not g159(n2068 ,n2067);
    not g160(n2066 ,n2065);
    not g161(n2064 ,n2063);
    not g162(n2062 ,n2061);
    not g163(n2060 ,n2059);
    nor g164(n2058 ,n674 ,n2041);
    nor g165(n2071 ,n698 ,n2038);
    nor g166(n2069 ,n871 ,n2037);
    nor g167(n2067 ,n672 ,n2036);
    nor g168(n2065 ,n805 ,n2039);
    nor g169(n2063 ,n873 ,n2040);
    nor g170(n2061 ,n828 ,n2035);
    nor g171(n2059 ,n744 ,n2026);
    not g172(n2057 ,n2056);
    not g173(n2055 ,n2054);
    not g174(n2053 ,n2052);
    not g175(n2051 ,n2050);
    not g176(n2049 ,n2048);
    not g177(n2047 ,n2046);
    not g178(n2045 ,n2044);
    not g179(n2043 ,n2042);
    nor g180(n2056 ,n801 ,n2029);
    nor g181(n2054 ,n833 ,n2032);
    nor g182(n2052 ,n705 ,n2031);
    nor g183(n2050 ,n794 ,n2030);
    nor g184(n2048 ,n810 ,n2033);
    nor g185(n2046 ,n907 ,n2028);
    nor g186(n2044 ,n837 ,n2027);
    nor g187(n2042 ,n663 ,n2034);
    or g188(n2041 ,n1752 ,n2019);
    or g189(n2040 ,n1755 ,n2020);
    or g190(n2039 ,n1770 ,n2017);
    or g191(n2038 ,n1767 ,n2024);
    or g192(n2037 ,n1764 ,n2023);
    or g193(n2036 ,n1761 ,n2022);
    or g194(n2035 ,n1758 ,n2021);
    or g195(n2034 ,n1724 ,n2010);
    or g196(n2033 ,n1746 ,n2025);
    or g197(n2032 ,n1743 ,n2008);
    or g198(n2031 ,n1739 ,n2015);
    or g199(n2030 ,n1736 ,n2014);
    or g200(n2029 ,n1733 ,n2013);
    or g201(n2028 ,n1730 ,n2012);
    or g202(n2027 ,n1727 ,n2011);
    or g203(n2026 ,n1749 ,n2018);
    or g204(n2025 ,n997 ,n2001);
    or g205(n2024 ,n1065 ,n1994);
    or g206(n2023 ,n1060 ,n1995);
    or g207(n2022 ,n1055 ,n1996);
    or g208(n2021 ,n1046 ,n1997);
    or g209(n2020 ,n1044 ,n1998);
    or g210(n2019 ,n1024 ,n1999);
    or g211(n2018 ,n1007 ,n2000);
    or g212(n2017 ,n1072 ,n1993);
    or g213(n2016 ,n1 ,n1991);
    or g214(n2015 ,n982 ,n2003);
    or g215(n2014 ,n975 ,n2004);
    or g216(n2013 ,n966 ,n2005);
    or g217(n2012 ,n961 ,n2006);
    or g218(n2011 ,n1011 ,n2007);
    or g219(n2010 ,n1079 ,n1992);
    nor g220(n2009 ,n1 ,n1990);
    or g221(n2008 ,n989 ,n2002);
    or g222(n2007 ,n669 ,n1973);
    or g223(n2006 ,n954 ,n1974);
    or g224(n2005 ,n816 ,n1975);
    or g225(n2004 ,n820 ,n1976);
    or g226(n2003 ,n904 ,n1977);
    or g227(n2002 ,n713 ,n1978);
    or g228(n2001 ,n722 ,n1979);
    or g229(n2000 ,n703 ,n1980);
    or g230(n1999 ,n848 ,n1981);
    or g231(n1998 ,n716 ,n1982);
    or g232(n1997 ,n925 ,n1983);
    or g233(n1996 ,n675 ,n1984);
    or g234(n1995 ,n921 ,n1985);
    or g235(n1994 ,n847 ,n1986);
    or g236(n1993 ,n943 ,n1987);
    or g237(n1992 ,n840 ,n1988);
    nor g238(n1991 ,n134 ,n1956);
    or g239(n1990 ,n134 ,n1972);
    or g240(n1989 ,n1430 ,n1475);
    or g241(n1988 ,n1772 ,n1771);
    or g242(n1987 ,n1769 ,n1768);
    or g243(n1986 ,n1766 ,n1765);
    or g244(n1985 ,n1763 ,n1762);
    or g245(n1984 ,n1760 ,n1759);
    or g246(n1983 ,n1757 ,n1756);
    or g247(n1982 ,n1754 ,n1753);
    or g248(n1981 ,n1751 ,n1750);
    or g249(n1980 ,n1748 ,n1747);
    or g250(n1979 ,n1745 ,n1744);
    or g251(n1978 ,n1741 ,n1740);
    or g252(n1977 ,n1738 ,n1737);
    or g253(n1976 ,n1735 ,n1734);
    or g254(n1975 ,n1732 ,n1731);
    or g255(n1974 ,n1729 ,n1728);
    or g256(n1973 ,n1726 ,n1725);
    or g257(n1972 ,n26[3] ,n1723);
    or g258(n1971 ,n1333 ,n1497);
    or g259(n1970 ,n1456 ,n1496);
    or g260(n1969 ,n1454 ,n1493);
    or g261(n1968 ,n1452 ,n1491);
    or g262(n1967 ,n651 ,n1488);
    or g263(n1966 ,n650 ,n1487);
    or g264(n1965 ,n645 ,n1485);
    or g265(n1964 ,n637 ,n1482);
    or g266(n1963 ,n638 ,n1481);
    or g267(n1962 ,n639 ,n1480);
    or g268(n1961 ,n643 ,n1479);
    or g269(n1960 ,n641 ,n1478);
    or g270(n1959 ,n644 ,n1477);
    or g271(n1958 ,n640 ,n1476);
    or g272(n1957 ,n1382 ,n1691);
    or g273(n1956 ,n26[3] ,n1742);
    or g274(n1955 ,n1419 ,n1717);
    or g275(n1954 ,n1428 ,n1720);
    or g276(n1953 ,n1425 ,n1719);
    or g277(n1952 ,n1426 ,n1718);
    or g278(n1951 ,n1424 ,n1716);
    or g279(n1950 ,n1421 ,n1714);
    or g280(n1949 ,n1423 ,n1715);
    or g281(n1948 ,n1417 ,n1713);
    or g282(n1947 ,n1413 ,n1712);
    or g283(n1946 ,n1411 ,n1710);
    or g284(n1945 ,n1412 ,n1711);
    or g285(n1944 ,n1409 ,n1709);
    or g286(n1943 ,n1408 ,n1707);
    or g287(n1942 ,n1406 ,n1705);
    or g288(n1941 ,n1407 ,n1708);
    or g289(n1940 ,n1427 ,n1704);
    or g290(n1939 ,n1405 ,n1706);
    or g291(n1938 ,n1404 ,n1702);
    or g292(n1937 ,n1403 ,n1703);
    or g293(n1936 ,n1173 ,n1701);
    or g294(n1935 ,n1400 ,n1700);
    or g295(n1934 ,n1398 ,n1699);
    or g296(n1933 ,n1397 ,n1582);
    or g297(n1932 ,n1395 ,n1780);
    or g298(n1931 ,n1393 ,n1697);
    or g299(n1930 ,n1379 ,n1692);
    or g300(n1929 ,n1385 ,n1695);
    or g301(n1928 ,n1384 ,n1694);
    or g302(n1927 ,n1383 ,n1693);
    or g303(n1926 ,n1381 ,n1689);
    or g304(n1925 ,n1270 ,n1777);
    or g305(n1924 ,n1378 ,n1688);
    or g306(n1923 ,n1377 ,n1686);
    or g307(n1922 ,n1376 ,n1687);
    or g308(n1921 ,n1373 ,n1683);
    or g309(n1920 ,n1375 ,n1685);
    or g310(n1919 ,n1374 ,n1684);
    or g311(n1918 ,n1372 ,n1681);
    or g312(n1917 ,n1370 ,n1680);
    or g313(n1916 ,n1371 ,n1682);
    or g314(n1915 ,n1368 ,n1679);
    or g315(n1914 ,n1364 ,n1678);
    or g316(n1913 ,n1361 ,n1677);
    or g317(n1912 ,n1360 ,n1676);
    or g318(n1911 ,n1357 ,n1675);
    or g319(n1910 ,n1358 ,n1674);
    or g320(n1909 ,n1356 ,n1673);
    or g321(n1908 ,n1353 ,n1671);
    or g322(n1907 ,n1354 ,n1672);
    or g323(n1906 ,n1352 ,n1670);
    or g324(n1905 ,n1350 ,n1668);
    or g325(n1904 ,n1351 ,n1669);
    or g326(n1903 ,n1348 ,n1667);
    or g327(n1902 ,n1347 ,n1666);
    or g328(n1901 ,n1346 ,n1665);
    or g329(n1900 ,n1343 ,n1664);
    or g330(n1899 ,n1341 ,n1663);
    or g331(n1898 ,n1330 ,n1662);
    or g332(n1897 ,n1322 ,n1655);
    or g333(n1896 ,n1327 ,n1659);
    or g334(n1895 ,n1328 ,n1661);
    or g335(n1894 ,n1326 ,n1660);
    or g336(n1893 ,n1325 ,n1658);
    or g337(n1892 ,n1324 ,n1657);
    or g338(n1891 ,n1323 ,n1656);
    or g339(n1890 ,n1320 ,n1653);
    or g340(n1889 ,n1321 ,n1654);
    or g341(n1888 ,n1319 ,n1652);
    or g342(n1887 ,n1318 ,n1648);
    or g343(n1886 ,n1317 ,n1651);
    or g344(n1885 ,n1316 ,n1650);
    or g345(n1884 ,n1315 ,n1649);
    or g346(n1883 ,n1311 ,n1643);
    or g347(n1882 ,n1313 ,n1645);
    or g348(n1881 ,n1314 ,n1647);
    or g349(n1880 ,n1312 ,n1646);
    or g350(n1879 ,n1309 ,n1644);
    or g351(n1878 ,n1304 ,n1638);
    or g352(n1877 ,n1305 ,n1642);
    or g353(n1876 ,n1302 ,n1641);
    or g354(n1875 ,n1300 ,n1640);
    or g355(n1874 ,n1294 ,n1635);
    or g356(n1873 ,n1298 ,n1637);
    or g357(n1872 ,n1299 ,n1639);
    or g358(n1871 ,n1297 ,n1636);
    or g359(n1870 ,n1295 ,n1632);
    or g360(n1869 ,n1296 ,n1634);
    or g361(n1868 ,n1279 ,n1626);
    or g362(n1867 ,n1293 ,n1633);
    or g363(n1866 ,n1291 ,n1630);
    or g364(n1865 ,n1292 ,n1631);
    or g365(n1864 ,n1289 ,n1628);
    or g366(n1863 ,n1290 ,n1629);
    or g367(n1862 ,n1288 ,n1627);
    or g368(n1861 ,n1286 ,n1625);
    or g369(n1860 ,n1283 ,n1773);
    or g370(n1859 ,n1285 ,n1624);
    or g371(n1858 ,n1282 ,n1698);
    or g372(n1857 ,n1276 ,n1774);
    or g373(n1856 ,n1273 ,n1775);
    or g374(n1855 ,n1271 ,n1776);
    or g375(n1854 ,n1269 ,n1541);
    or g376(n1853 ,n1380 ,n1690);
    or g377(n1852 ,n1266 ,n1778);
    or g378(n1851 ,n1268 ,n1779);
    or g379(n1850 ,n1267 ,n1622);
    or g380(n1849 ,n1265 ,n1619);
    or g381(n1848 ,n1264 ,n1621);
    or g382(n1847 ,n1262 ,n1617);
    or g383(n1846 ,n1263 ,n1618);
    or g384(n1845 ,n1261 ,n1616);
    or g385(n1844 ,n1259 ,n1615);
    or g386(n1843 ,n1255 ,n1610);
    or g387(n1842 ,n1258 ,n1614);
    or g388(n1841 ,n1257 ,n1613);
    or g389(n1840 ,n1254 ,n1611);
    or g390(n1839 ,n1256 ,n1612);
    or g391(n1838 ,n1260 ,n1620);
    or g392(n1837 ,n1252 ,n1609);
    or g393(n1836 ,n1250 ,n1607);
    or g394(n1835 ,n1248 ,n1606);
    or g395(n1834 ,n1246 ,n1605);
    or g396(n1833 ,n1245 ,n1604);
    or g397(n1832 ,n1243 ,n1603);
    or g398(n1831 ,n1244 ,n1608);
    or g399(n1830 ,n1238 ,n1601);
    or g400(n1829 ,n1236 ,n1602);
    or g401(n1828 ,n1234 ,n1600);
    or g402(n1827 ,n1235 ,n1599);
    or g403(n1826 ,n1224 ,n1589);
    or g404(n1825 ,n1396 ,n1598);
    or g405(n1824 ,n1233 ,n1596);
    or g406(n1823 ,n1232 ,n1595);
    or g407(n1822 ,n1231 ,n1594);
    or g408(n1821 ,n1229 ,n1592);
    or g409(n1820 ,n1230 ,n1593);
    or g410(n1819 ,n1228 ,n1591);
    or g411(n1818 ,n1227 ,n1587);
    or g412(n1817 ,n1226 ,n1590);
    or g413(n1816 ,n1225 ,n1588);
    or g414(n1815 ,n1223 ,n1586);
    or g415(n1814 ,n1221 ,n1585);
    or g416(n1813 ,n1222 ,n1584);
    or g417(n1812 ,n1217 ,n1581);
    or g418(n1811 ,n1219 ,n1583);
    or g419(n1810 ,n1214 ,n1580);
    or g420(n1809 ,n1213 ,n1578);
    or g421(n1808 ,n1209 ,n1576);
    or g422(n1807 ,n1211 ,n1579);
    or g423(n1806 ,n1210 ,n1577);
    or g424(n1805 ,n1197 ,n1575);
    or g425(n1804 ,n1196 ,n1574);
    or g426(n1803 ,n1195 ,n1573);
    or g427(n1802 ,n1193 ,n1570);
    or g428(n1801 ,n1194 ,n1572);
    or g429(n1800 ,n1192 ,n1571);
    or g430(n1799 ,n1191 ,n1569);
    or g431(n1798 ,n1189 ,n1568);
    or g432(n1797 ,n1187 ,n1563);
    or g433(n1796 ,n1188 ,n1567);
    or g434(n1795 ,n1185 ,n1566);
    or g435(n1794 ,n1184 ,n1565);
    or g436(n1793 ,n1169 ,n1561);
    or g437(n1792 ,n1174 ,n1562);
    or g438(n1791 ,n1171 ,n1559);
    or g439(n1790 ,n1168 ,n1557);
    or g440(n1789 ,n1175 ,n1560);
    or g441(n1788 ,n1164 ,n1564);
    or g442(n1787 ,n1167 ,n1558);
    or g443(n1786 ,n1165 ,n1554);
    or g444(n1785 ,n1166 ,n1556);
    or g445(n1784 ,n1163 ,n1555);
    or g446(n1783 ,n1172 ,n1696);
    or g447(n1782 ,n1249 ,n1721);
    or g448(n1781 ,n1162 ,n1597);
    nor g449(n1780 ,n776 ,n1200);
    nor g450(n1779 ,n778 ,n1206);
    nor g451(n1778 ,n760 ,n1198);
    nor g452(n1777 ,n778 ,n1208);
    nor g453(n1776 ,n778 ,n1202);
    nor g454(n1775 ,n778 ,n1205);
    nor g455(n1774 ,n760 ,n1199);
    nor g456(n1773 ,n760 ,n1204);
    or g457(n1772 ,n1047 ,n1078);
    or g458(n1771 ,n960 ,n1077);
    or g459(n1770 ,n1022 ,n1073);
    or g460(n1769 ,n1027 ,n1071);
    or g461(n1768 ,n1028 ,n1029);
    or g462(n1767 ,n1067 ,n1066);
    or g463(n1766 ,n1039 ,n1032);
    or g464(n1765 ,n1033 ,n1062);
    or g465(n1764 ,n1036 ,n1040);
    or g466(n1763 ,n1051 ,n1056);
    or g467(n1762 ,n1059 ,n1058);
    or g468(n1761 ,n992 ,n1075);
    or g469(n1760 ,n1070 ,n970);
    or g470(n1759 ,n1054 ,n1053);
    or g471(n1758 ,n1050 ,n1048);
    or g472(n1757 ,n1068 ,n1052);
    or g473(n1756 ,n990 ,n1045);
    or g474(n1755 ,n977 ,n1035);
    or g475(n1754 ,n983 ,n969);
    or g476(n1753 ,n1043 ,n1042);
    or g477(n1752 ,n1000 ,n968);
    or g478(n1751 ,n1057 ,n1038);
    or g479(n1750 ,n1037 ,n1069);
    or g480(n1749 ,n1010 ,n1009);
    or g481(n1748 ,n1005 ,n1004);
    or g482(n1747 ,n1003 ,n1002);
    or g483(n1746 ,n999 ,n998);
    or g484(n1745 ,n1064 ,n996);
    or g485(n1744 ,n995 ,n994);
    or g486(n1743 ,n991 ,n1031);
    or g487(n1742 ,n600 ,n1144);
    or g488(n1741 ,n988 ,n987);
    or g489(n1740 ,n986 ,n985);
    or g490(n1739 ,n1041 ,n1023);
    or g491(n1738 ,n981 ,n980);
    or g492(n1737 ,n979 ,n978);
    or g493(n1736 ,n993 ,n1012);
    or g494(n1735 ,n974 ,n973);
    or g495(n1734 ,n972 ,n971);
    or g496(n1733 ,n1014 ,n967);
    or g497(n1732 ,n965 ,n1026);
    or g498(n1731 ,n964 ,n963);
    or g499(n1730 ,n1063 ,n1034);
    or g500(n1729 ,n1049 ,n959);
    or g501(n1728 ,n1074 ,n958);
    or g502(n1727 ,n1001 ,n962);
    or g503(n1726 ,n984 ,n1017);
    or g504(n1725 ,n976 ,n1025);
    or g505(n1724 ,n1006 ,n1008);
    or g506(n1723 ,n26[0] ,n1161);
    nor g507(n1722 ,n1 ,n1076);
    nor g508(n1721 ,n752 ,n1206);
    nor g509(n1720 ,n766 ,n1199);
    nor g510(n1719 ,n766 ,n1198);
    nor g511(n1718 ,n752 ,n1207);
    nor g512(n1717 ,n780 ,n1199);
    nor g513(n1716 ,n766 ,n1201);
    nor g514(n1715 ,n766 ,n1200);
    nor g515(n1714 ,n752 ,n1203);
    nor g516(n1713 ,n752 ,n1204);
    nor g517(n1712 ,n752 ,n1199);
    nor g518(n1711 ,n752 ,n1198);
    nor g519(n1710 ,n776 ,n1205);
    nor g520(n1709 ,n776 ,n1202);
    nor g521(n1708 ,n776 ,n1208);
    nor g522(n1707 ,n780 ,n1198);
    nor g523(n1706 ,n776 ,n1206);
    nor g524(n1705 ,n752 ,n1201);
    nor g525(n1704 ,n776 ,n1207);
    nor g526(n1703 ,n776 ,n1203);
    nor g527(n1702 ,n752 ,n1200);
    nor g528(n1701 ,n776 ,n1204);
    nor g529(n1700 ,n776 ,n1199);
    nor g530(n1699 ,n776 ,n1198);
    nor g531(n1698 ,n764 ,n1200);
    nor g532(n1697 ,n780 ,n1201);
    nor g533(n1696 ,n754 ,n1205);
    nor g534(n1695 ,n754 ,n1202);
    nor g535(n1694 ,n750 ,n1205);
    nor g536(n1693 ,n754 ,n1208);
    nor g537(n1692 ,n780 ,n1200);
    nor g538(n1691 ,n754 ,n1206);
    nor g539(n1690 ,n754 ,n1207);
    nor g540(n1689 ,n750 ,n1202);
    nor g541(n1688 ,n754 ,n1203);
    nor g542(n1687 ,n754 ,n1204);
    nor g543(n1686 ,n750 ,n1208);
    nor g544(n1685 ,n754 ,n1199);
    nor g545(n1684 ,n754 ,n1198);
    nor g546(n1683 ,n750 ,n1206);
    nor g547(n1682 ,n750 ,n1207);
    nor g548(n1681 ,n754 ,n1201);
    nor g549(n1680 ,n754 ,n1200);
    nor g550(n1679 ,n750 ,n1203);
    nor g551(n1678 ,n750 ,n1204);
    nor g552(n1677 ,n750 ,n1199);
    nor g553(n1676 ,n758 ,n1205);
    nor g554(n1675 ,n758 ,n1202);
    nor g555(n1674 ,n750 ,n1198);
    nor g556(n1673 ,n758 ,n1208);
    nor g557(n1672 ,n758 ,n1206);
    nor g558(n1671 ,n750 ,n1201);
    nor g559(n1670 ,n758 ,n1207);
    nor g560(n1669 ,n758 ,n1203);
    nor g561(n1668 ,n750 ,n1200);
    nor g562(n1667 ,n758 ,n1204);
    nor g563(n1666 ,n758 ,n1199);
    nor g564(n1665 ,n758 ,n1198);
    nor g565(n1664 ,n758 ,n1201);
    nor g566(n1663 ,n758 ,n1200);
    nor g567(n1662 ,n756 ,n1205);
    nor g568(n1661 ,n756 ,n1202);
    nor g569(n1660 ,n756 ,n1208);
    nor g570(n1659 ,n762 ,n1205);
    nor g571(n1658 ,n756 ,n1206);
    nor g572(n1657 ,n762 ,n1202);
    nor g573(n1656 ,n756 ,n1207);
    nor g574(n1655 ,n760 ,n1205);
    nor g575(n1654 ,n756 ,n1203);
    nor g576(n1653 ,n762 ,n1208);
    nor g577(n1652 ,n756 ,n1204);
    nor g578(n1651 ,n756 ,n1199);
    nor g579(n1650 ,n762 ,n1206);
    nor g580(n1649 ,n756 ,n1198);
    nor g581(n1648 ,n760 ,n1202);
    nor g582(n1647 ,n756 ,n1201);
    nor g583(n1646 ,n756 ,n1200);
    nor g584(n1645 ,n762 ,n1207);
    nor g585(n1644 ,n762 ,n1203);
    nor g586(n1643 ,n760 ,n1208);
    nor g587(n1642 ,n762 ,n1204);
    nor g588(n1641 ,n762 ,n1199);
    nor g589(n1640 ,n764 ,n1205);
    nor g590(n1639 ,n764 ,n1202);
    nor g591(n1638 ,n760 ,n1206);
    nor g592(n1637 ,n762 ,n1198);
    nor g593(n1636 ,n764 ,n1208);
    nor g594(n1635 ,n760 ,n1207);
    nor g595(n1634 ,n764 ,n1206);
    nor g596(n1633 ,n764 ,n1207);
    nor g597(n1632 ,n762 ,n1201);
    nor g598(n1631 ,n764 ,n1203);
    nor g599(n1630 ,n762 ,n1200);
    nor g600(n1629 ,n764 ,n1204);
    nor g601(n1628 ,n760 ,n1203);
    nor g602(n1627 ,n764 ,n1199);
    nor g603(n1626 ,n780 ,n1205);
    nor g604(n1625 ,n764 ,n1198);
    nor g605(n1624 ,n764 ,n1201);
    or g606(n1623 ,n1388 ,n1133);
    nor g607(n1622 ,n778 ,n1207);
    nor g608(n1621 ,n778 ,n1203);
    nor g609(n1620 ,n760 ,n1201);
    nor g610(n1619 ,n770 ,n1202);
    nor g611(n1618 ,n778 ,n1204);
    nor g612(n1617 ,n770 ,n1208);
    nor g613(n1616 ,n778 ,n1199);
    nor g614(n1615 ,n778 ,n1198);
    nor g615(n1614 ,n770 ,n1206);
    nor g616(n1613 ,n778 ,n1201);
    nor g617(n1612 ,n778 ,n1200);
    nor g618(n1611 ,n770 ,n1207);
    nor g619(n1610 ,n760 ,n1200);
    nor g620(n1609 ,n770 ,n1203);
    nor g621(n1608 ,n780 ,n1202);
    nor g622(n1607 ,n770 ,n1204);
    nor g623(n1606 ,n770 ,n1199);
    nor g624(n1605 ,n770 ,n1198);
    nor g625(n1604 ,n770 ,n1201);
    nor g626(n1603 ,n770 ,n1200);
    nor g627(n1602 ,n772 ,n1205);
    nor g628(n1601 ,n780 ,n1208);
    nor g629(n1600 ,n774 ,n1205);
    nor g630(n1599 ,n772 ,n1202);
    nor g631(n1598 ,n772 ,n1208);
    nor g632(n1597 ,n766 ,n1204);
    nor g633(n1596 ,n774 ,n1202);
    nor g634(n1595 ,n772 ,n1206);
    nor g635(n1594 ,n772 ,n1207);
    nor g636(n1593 ,n772 ,n1203);
    nor g637(n1592 ,n774 ,n1208);
    nor g638(n1591 ,n772 ,n1204);
    nor g639(n1590 ,n772 ,n1199);
    nor g640(n1589 ,n780 ,n1206);
    nor g641(n1588 ,n772 ,n1198);
    nor g642(n1587 ,n774 ,n1206);
    nor g643(n1586 ,n772 ,n1201);
    nor g644(n1585 ,n774 ,n1207);
    nor g645(n1584 ,n772 ,n1200);
    nor g646(n1583 ,n774 ,n1203);
    nor g647(n1582 ,n776 ,n1201);
    nor g648(n1581 ,n774 ,n1204);
    nor g649(n1580 ,n774 ,n1199);
    nor g650(n1579 ,n768 ,n1205);
    nor g651(n1578 ,n780 ,n1207);
    nor g652(n1577 ,n768 ,n1202);
    nor g653(n1576 ,n774 ,n1198);
    nor g654(n1575 ,n768 ,n1208);
    nor g655(n1574 ,n774 ,n1201);
    nor g656(n1573 ,n768 ,n1206);
    nor g657(n1572 ,n768 ,n1207);
    nor g658(n1571 ,n768 ,n1203);
    nor g659(n1570 ,n774 ,n1200);
    nor g660(n1569 ,n768 ,n1204);
    nor g661(n1568 ,n768 ,n1199);
    nor g662(n1567 ,n768 ,n1198);
    nor g663(n1566 ,n768 ,n1201);
    nor g664(n1565 ,n768 ,n1200);
    nor g665(n1564 ,n766 ,n1208);
    nor g666(n1563 ,n780 ,n1203);
    nor g667(n1562 ,n766 ,n1205);
    nor g668(n1561 ,n780 ,n1204);
    nor g669(n1560 ,n752 ,n1205);
    nor g670(n1559 ,n766 ,n1202);
    nor g671(n1558 ,n766 ,n1206);
    nor g672(n1557 ,n752 ,n1202);
    nor g673(n1556 ,n766 ,n1207);
    nor g674(n1555 ,n766 ,n1203);
    nor g675(n1554 ,n752 ,n1208);
    or g676(n1553 ,n1420 ,n1160);
    or g677(n1552 ,n1418 ,n1143);
    or g678(n1551 ,n1416 ,n1142);
    or g679(n1550 ,n1415 ,n1141);
    or g680(n1549 ,n1414 ,n1140);
    or g681(n1548 ,n1401 ,n1159);
    or g682(n1547 ,n1399 ,n1087);
    or g683(n1546 ,n1394 ,n1158);
    or g684(n1545 ,n1392 ,n1135);
    or g685(n1544 ,n1391 ,n1137);
    or g686(n1543 ,n1389 ,n1134);
    or g687(n1542 ,n1410 ,n1131);
    nor g688(n1541 ,n770 ,n1205);
    or g689(n1540 ,n1386 ,n1089);
    or g690(n1539 ,n1387 ,n1132);
    or g691(n1538 ,n1366 ,n1155);
    or g692(n1537 ,n1369 ,n1156);
    or g693(n1536 ,n1367 ,n1130);
    or g694(n1535 ,n1355 ,n1124);
    or g695(n1534 ,n1365 ,n1129);
    or g696(n1533 ,n1363 ,n1128);
    or g697(n1532 ,n1362 ,n1126);
    or g698(n1531 ,n1359 ,n1125);
    or g699(n1530 ,n1349 ,n1123);
    or g700(n1529 ,n1345 ,n1154);
    or g701(n1528 ,n1344 ,n1122);
    or g702(n1527 ,n1339 ,n1153);
    or g703(n1526 ,n1338 ,n1121);
    or g704(n1525 ,n1337 ,n1120);
    or g705(n1524 ,n1340 ,n1119);
    or g706(n1523 ,n1335 ,n1117);
    or g707(n1522 ,n1336 ,n1118);
    or g708(n1521 ,n1334 ,n1138);
    or g709(n1520 ,n1458 ,n1113);
    or g710(n1519 ,n1332 ,n1116);
    or g711(n1518 ,n1331 ,n1115);
    or g712(n1517 ,n1342 ,n1114);
    or g713(n1516 ,n1308 ,n1109);
    or g714(n1515 ,n1310 ,n1146);
    or g715(n1514 ,n1307 ,n1112);
    or g716(n1513 ,n1306 ,n1111);
    or g717(n1512 ,n1303 ,n1110);
    or g718(n1511 ,n1301 ,n1108);
    or g719(n1510 ,n1287 ,n1152);
    or g720(n1509 ,n1284 ,n1107);
    or g721(n1508 ,n1281 ,n1151);
    or g722(n1507 ,n1280 ,n1084);
    or g723(n1506 ,n1278 ,n1106);
    or g724(n1505 ,n1277 ,n1105);
    or g725(n1504 ,n1170 ,n1104);
    or g726(n1503 ,n1274 ,n1102);
    or g727(n1502 ,n1275 ,n1103);
    or g728(n1501 ,n1272 ,n1101);
    or g729(n1500 ,n1253 ,n1150);
    or g730(n1499 ,n1251 ,n1149);
    or g731(n1498 ,n1247 ,n1100);
    or g732(n1497 ,n646 ,n1457);
    or g733(n1496 ,n647 ,n1455);
    or g734(n1495 ,n1241 ,n1148);
    or g735(n1494 ,n1402 ,n1098);
    or g736(n1493 ,n642 ,n1453);
    or g737(n1492 ,n1242 ,n1099);
    or g738(n1491 ,n649 ,n1451);
    or g739(n1490 ,n1240 ,n1097);
    or g740(n1489 ,n1239 ,n1096);
    or g741(n1488 ,n1450 ,n1449);
    or g742(n1487 ,n1447 ,n1448);
    or g743(n1486 ,n1422 ,n1092);
    or g744(n1485 ,n1446 ,n1445);
    or g745(n1484 ,n1180 ,n1095);
    or g746(n1483 ,n1237 ,n1088);
    or g747(n1482 ,n1443 ,n1444);
    or g748(n1481 ,n1442 ,n1441);
    or g749(n1480 ,n1440 ,n1439);
    or g750(n1479 ,n1438 ,n1437);
    or g751(n1478 ,n1436 ,n1435);
    or g752(n1477 ,n1434 ,n1433);
    or g753(n1476 ,n1432 ,n1431);
    or g754(n1475 ,n648 ,n1429);
    or g755(n1474 ,n1390 ,n1127);
    or g756(n1473 ,n1220 ,n1147);
    or g757(n1472 ,n1218 ,n1094);
    or g758(n1471 ,n1216 ,n1093);
    or g759(n1470 ,n1215 ,n1091);
    or g760(n1469 ,n1212 ,n1090);
    or g761(n1468 ,n1190 ,n1157);
    or g762(n1467 ,n1186 ,n1086);
    or g763(n1466 ,n1183 ,n1085);
    or g764(n1465 ,n1329 ,n1145);
    or g765(n1464 ,n1182 ,n1083);
    or g766(n1463 ,n1181 ,n1081);
    or g767(n1462 ,n1176 ,n1080);
    or g768(n1461 ,n1179 ,n1082);
    or g769(n1460 ,n1178 ,n1139);
    or g770(n1459 ,n1177 ,n1136);
    nor g771(n1458 ,n214 ,n761);
    nor g772(n1457 ,n292 ,n787);
    nor g773(n1456 ,n286 ,n787);
    nor g774(n1455 ,n320 ,n786);
    nor g775(n1454 ,n283 ,n787);
    nor g776(n1453 ,n319 ,n786);
    nor g777(n1452 ,n297 ,n787);
    nor g778(n1451 ,n152 ,n786);
    nor g779(n1450 ,n327 ,n786);
    nor g780(n1449 ,n302 ,n787);
    nor g781(n1448 ,n280 ,n787);
    nor g782(n1447 ,n324 ,n786);
    nor g783(n1446 ,n169 ,n786);
    nor g784(n1445 ,n296 ,n787);
    nor g785(n1444 ,n312 ,n787);
    nor g786(n1443 ,n326 ,n786);
    nor g787(n1442 ,n172 ,n786);
    nor g788(n1441 ,n282 ,n787);
    nor g789(n1440 ,n171 ,n786);
    nor g790(n1439 ,n284 ,n787);
    nor g791(n1438 ,n325 ,n786);
    nor g792(n1437 ,n313 ,n787);
    nor g793(n1436 ,n167 ,n786);
    nor g794(n1435 ,n307 ,n787);
    nor g795(n1434 ,n323 ,n786);
    nor g796(n1433 ,n289 ,n787);
    nor g797(n1432 ,n322 ,n786);
    nor g798(n1431 ,n299 ,n787);
    nor g799(n1430 ,n314 ,n787);
    nor g800(n1429 ,n160 ,n786);
    nor g801(n1428 ,n223 ,n767);
    nor g802(n1427 ,n275 ,n777);
    nor g803(n1426 ,n345 ,n753);
    nor g804(n1425 ,n256 ,n767);
    nor g805(n1424 ,n442 ,n767);
    nor g806(n1423 ,n374 ,n767);
    nor g807(n1422 ,n428 ,n773);
    nor g808(n1421 ,n276 ,n753);
    nor g809(n1420 ,n393 ,n767);
    nor g810(n1419 ,n479 ,n781);
    nor g811(n1418 ,n371 ,n777);
    nor g812(n1417 ,n178 ,n753);
    nor g813(n1416 ,n201 ,n777);
    nor g814(n1415 ,n350 ,n777);
    nor g815(n1414 ,n173 ,n777);
    nor g816(n1413 ,n401 ,n753);
    nor g817(n1412 ,n490 ,n753);
    nor g818(n1411 ,n340 ,n777);
    nor g819(n1410 ,n358 ,n751);
    nor g820(n1409 ,n448 ,n777);
    nor g821(n1408 ,n363 ,n781);
    nor g822(n1407 ,n238 ,n777);
    nor g823(n1406 ,n334 ,n753);
    nor g824(n1405 ,n215 ,n777);
    nor g825(n1404 ,n251 ,n753);
    nor g826(n1403 ,n414 ,n777);
    nor g827(n1402 ,n186 ,n773);
    nor g828(n1401 ,n226 ,n753);
    nor g829(n1400 ,n220 ,n777);
    nor g830(n1399 ,n485 ,n751);
    nor g831(n1398 ,n406 ,n777);
    nor g832(n1397 ,n356 ,n777);
    nor g833(n1396 ,n174 ,n773);
    nor g834(n1395 ,n189 ,n777);
    nor g835(n1394 ,n349 ,n777);
    nor g836(n1393 ,n388 ,n781);
    nor g837(n1392 ,n402 ,n751);
    nor g838(n1391 ,n404 ,n755);
    nor g839(n1390 ,n208 ,n781);
    nor g840(n1389 ,n343 ,n755);
    nor g841(n1388 ,n332 ,n755);
    nor g842(n1387 ,n369 ,n755);
    nor g843(n1386 ,n494 ,n751);
    nor g844(n1385 ,n183 ,n755);
    nor g845(n1384 ,n434 ,n751);
    nor g846(n1383 ,n269 ,n755);
    nor g847(n1382 ,n203 ,n755);
    nor g848(n1381 ,n489 ,n751);
    nor g849(n1380 ,n468 ,n755);
    nor g850(n1379 ,n471 ,n781);
    nor g851(n1378 ,n445 ,n755);
    nor g852(n1377 ,n209 ,n751);
    nor g853(n1376 ,n192 ,n755);
    nor g854(n1375 ,n493 ,n755);
    nor g855(n1374 ,n502 ,n755);
    nor g856(n1373 ,n486 ,n751);
    nor g857(n1372 ,n235 ,n755);
    nor g858(n1371 ,n423 ,n751);
    nor g859(n1370 ,n175 ,n755);
    nor g860(n1369 ,n330 ,n755);
    nor g861(n1368 ,n216 ,n751);
    nor g862(n1367 ,n331 ,n759);
    nor g863(n1366 ,n338 ,n781);
    nor g864(n1365 ,n263 ,n759);
    nor g865(n1364 ,n274 ,n751);
    nor g866(n1363 ,n191 ,n759);
    nor g867(n1362 ,n458 ,n759);
    nor g868(n1361 ,n378 ,n751);
    nor g869(n1360 ,n480 ,n759);
    nor g870(n1359 ,n386 ,n761);
    nor g871(n1358 ,n243 ,n751);
    nor g872(n1357 ,n491 ,n759);
    nor g873(n1356 ,n242 ,n759);
    nor g874(n1355 ,n437 ,n781);
    nor g875(n1354 ,n333 ,n759);
    nor g876(n1353 ,n368 ,n751);
    nor g877(n1352 ,n341 ,n759);
    nor g878(n1351 ,n384 ,n759);
    nor g879(n1350 ,n373 ,n751);
    nor g880(n1349 ,n377 ,n761);
    nor g881(n1348 ,n447 ,n759);
    nor g882(n1347 ,n197 ,n759);
    nor g883(n1346 ,n412 ,n759);
    nor g884(n1345 ,n357 ,n751);
    nor g885(n1344 ,n194 ,n763);
    nor g886(n1343 ,n488 ,n759);
    nor g887(n1342 ,n206 ,n781);
    nor g888(n1341 ,n415 ,n759);
    nor g889(n1340 ,n483 ,n761);
    nor g890(n1339 ,n459 ,n759);
    nor g891(n1338 ,n424 ,n763);
    nor g892(n1337 ,n400 ,n757);
    nor g893(n1336 ,n277 ,n757);
    nor g894(n1335 ,n176 ,n763);
    nor g895(n1334 ,n237 ,n757);
    nor g896(n1333 ,n321 ,n786);
    nor g897(n1332 ,n245 ,n757);
    nor g898(n1331 ,n451 ,n763);
    nor g899(n1330 ,n430 ,n757);
    nor g900(n1329 ,n267 ,n769);
    nor g901(n1328 ,n181 ,n757);
    nor g902(n1327 ,n367 ,n763);
    nor g903(n1326 ,n409 ,n757);
    nor g904(n1325 ,n359 ,n757);
    nor g905(n1324 ,n264 ,n763);
    nor g906(n1323 ,n433 ,n757);
    nor g907(n1322 ,n441 ,n761);
    nor g908(n1321 ,n443 ,n757);
    nor g909(n1320 ,n328 ,n763);
    nor g910(n1319 ,n255 ,n757);
    nor g911(n1318 ,n461 ,n761);
    nor g912(n1317 ,n422 ,n757);
    nor g913(n1316 ,n339 ,n763);
    nor g914(n1315 ,n405 ,n757);
    nor g915(n1314 ,n410 ,n757);
    nor g916(n1313 ,n417 ,n763);
    nor g917(n1312 ,n481 ,n757);
    nor g918(n1311 ,n407 ,n761);
    nor g919(n1310 ,n469 ,n757);
    nor g920(n1309 ,n413 ,n763);
    nor g921(n1308 ,n249 ,n781);
    nor g922(n1307 ,n212 ,n765);
    nor g923(n1306 ,n195 ,n765);
    nor g924(n1305 ,n262 ,n763);
    nor g925(n1304 ,n432 ,n761);
    nor g926(n1303 ,n429 ,n765);
    nor g927(n1302 ,n248 ,n763);
    nor g928(n1301 ,n180 ,n765);
    nor g929(n1300 ,n416 ,n765);
    nor g930(n1299 ,n403 ,n765);
    nor g931(n1298 ,n501 ,n763);
    nor g932(n1297 ,n348 ,n765);
    nor g933(n1296 ,n184 ,n765);
    nor g934(n1295 ,n360 ,n763);
    nor g935(n1294 ,n498 ,n761);
    nor g936(n1293 ,n342 ,n765);
    nor g937(n1292 ,n390 ,n765);
    nor g938(n1291 ,n499 ,n763);
    nor g939(n1290 ,n354 ,n765);
    nor g940(n1289 ,n453 ,n761);
    nor g941(n1288 ,n450 ,n765);
    nor g942(n1287 ,n265 ,n763);
    nor g943(n1286 ,n439 ,n765);
    nor g944(n1285 ,n207 ,n765);
    nor g945(n1284 ,n347 ,n771);
    nor g946(n1283 ,n224 ,n761);
    nor g947(n1282 ,n456 ,n765);
    nor g948(n1281 ,n362 ,n765);
    nor g949(n1280 ,n257 ,n779);
    nor g950(n1279 ,n478 ,n781);
    nor g951(n1278 ,n457 ,n771);
    nor g952(n1277 ,n222 ,n779);
    nor g953(n1276 ,n376 ,n761);
    nor g954(n1275 ,n177 ,n779);
    nor g955(n1274 ,n392 ,n771);
    nor g956(n1273 ,n351 ,n779);
    nor g957(n1272 ,n221 ,n771);
    nor g958(n1271 ,n266 ,n779);
    nor g959(n1270 ,n205 ,n779);
    nor g960(n1269 ,n253 ,n771);
    nor g961(n1268 ,n185 ,n779);
    nor g962(n1267 ,n455 ,n779);
    nor g963(n1266 ,n366 ,n761);
    nor g964(n1265 ,n202 ,n771);
    nor g965(n1264 ,n463 ,n779);
    nor g966(n1263 ,n419 ,n779);
    nor g967(n1262 ,n408 ,n771);
    nor g968(n1261 ,n380 ,n779);
    nor g969(n1260 ,n492 ,n761);
    nor g970(n1259 ,n438 ,n779);
    nor g971(n1258 ,n268 ,n771);
    nor g972(n1257 ,n250 ,n779);
    nor g973(n1256 ,n239 ,n779);
    nor g974(n1255 ,n464 ,n761);
    nor g975(n1254 ,n187 ,n771);
    nor g976(n1253 ,n225 ,n779);
    nor g977(n1252 ,n381 ,n771);
    nor g978(n1251 ,n329 ,n761);
    nor g979(n1250 ,n336 ,n771);
    nor g980(n1249 ,n440 ,n753);
    nor g981(n1248 ,n444 ,n771);
    nor g982(n1247 ,n241 ,n775);
    nor g983(n1246 ,n396 ,n771);
    nor g984(n1245 ,n372 ,n771);
    nor g985(n1244 ,n411 ,n781);
    nor g986(n1243 ,n353 ,n771);
    nor g987(n1242 ,n272 ,n775);
    nor g988(n1241 ,n199 ,n771);
    nor g989(n1240 ,n382 ,n773);
    nor g990(n1239 ,n462 ,n775);
    nor g991(n1238 ,n467 ,n781);
    nor g992(n1237 ,n446 ,n773);
    nor g993(n1236 ,n364 ,n773);
    nor g994(n1235 ,n211 ,n773);
    nor g995(n1234 ,n395 ,n775);
    nor g996(n1233 ,n190 ,n775);
    nor g997(n1232 ,n425 ,n773);
    nor g998(n1231 ,n227 ,n773);
    nor g999(n1230 ,n427 ,n773);
    nor g1000(n1229 ,n431 ,n775);
    nor g1001(n1228 ,n418 ,n773);
    nor g1002(n1227 ,n476 ,n775);
    nor g1003(n1226 ,n182 ,n773);
    nor g1004(n1225 ,n335 ,n773);
    nor g1005(n1224 ,n229 ,n781);
    nor g1006(n1223 ,n398 ,n773);
    nor g1007(n1222 ,n244 ,n773);
    nor g1008(n1221 ,n497 ,n775);
    nor g1009(n1220 ,n466 ,n773);
    nor g1010(n1219 ,n231 ,n775);
    nor g1011(n1218 ,n477 ,n769);
    nor g1012(n1217 ,n420 ,n775);
    nor g1013(n1216 ,n232 ,n769);
    nor g1014(n1215 ,n397 ,n769);
    nor g1015(n1214 ,n365 ,n775);
    nor g1016(n1213 ,n474 ,n781);
    nor g1017(n1212 ,n387 ,n769);
    nor g1018(n1211 ,n436 ,n769);
    nor g1019(n1210 ,n394 ,n769);
    nor g1020(n1209 ,n188 ,n775);
    nor g1021(n1197 ,n240 ,n769);
    nor g1022(n1196 ,n204 ,n775);
    nor g1023(n1195 ,n200 ,n769);
    nor g1024(n1194 ,n465 ,n769);
    nor g1025(n1193 ,n352 ,n775);
    nor g1026(n1192 ,n219 ,n769);
    nor g1027(n1191 ,n230 ,n769);
    nor g1028(n1190 ,n399 ,n775);
    nor g1029(n1189 ,n472 ,n769);
    nor g1030(n1188 ,n273 ,n769);
    nor g1031(n1187 ,n234 ,n781);
    nor g1032(n1186 ,n475 ,n753);
    nor g1033(n1185 ,n449 ,n769);
    nor g1034(n1184 ,n228 ,n769);
    nor g1035(n1183 ,n246 ,n753);
    nor g1036(n1182 ,n454 ,n767);
    nor g1037(n1181 ,n271 ,n753);
    nor g1038(n1180 ,n500 ,n775);
    nor g1039(n1179 ,n421 ,n767);
    nor g1040(n1178 ,n452 ,n767);
    nor g1041(n1177 ,n496 ,n767);
    nor g1042(n1176 ,n259 ,n753);
    nor g1043(n1175 ,n247 ,n753);
    nor g1044(n1174 ,n260 ,n767);
    nor g1045(n1173 ,n385 ,n777);
    nor g1046(n1172 ,n270 ,n755);
    nor g1047(n1171 ,n236 ,n767);
    nor g1048(n1170 ,n379 ,n779);
    nor g1049(n1169 ,n355 ,n781);
    nor g1050(n1168 ,n213 ,n753);
    nor g1051(n1167 ,n375 ,n767);
    nor g1052(n1166 ,n435 ,n767);
    nor g1053(n1165 ,n391 ,n753);
    nor g1054(n1164 ,n196 ,n767);
    nor g1055(n1163 ,n487 ,n767);
    nor g1056(n1162 ,n473 ,n767);
    or g1057(n1161 ,n788 ,n618);
    nor g1058(n1160 ,n135 ,n766);
    nor g1059(n1159 ,n135 ,n752);
    nor g1060(n1158 ,n135 ,n776);
    nor g1061(n1157 ,n135 ,n774);
    nor g1062(n1156 ,n135 ,n754);
    nor g1063(n1155 ,n135 ,n780);
    nor g1064(n1154 ,n135 ,n750);
    nor g1065(n1153 ,n135 ,n758);
    nor g1066(n1152 ,n135 ,n762);
    nor g1067(n1151 ,n135 ,n764);
    nor g1068(n1150 ,n135 ,n778);
    nor g1069(n1149 ,n135 ,n760);
    nor g1070(n1148 ,n135 ,n770);
    nor g1071(n1147 ,n135 ,n772);
    nor g1072(n1146 ,n135 ,n756);
    nor g1073(n1145 ,n135 ,n768);
    or g1074(n1144 ,n26[4] ,n606);
    nor g1075(n1143 ,n564 ,n776);
    nor g1076(n1142 ,n567 ,n776);
    nor g1077(n1141 ,n566 ,n776);
    nor g1078(n1140 ,n565 ,n776);
    nor g1079(n1139 ,n566 ,n766);
    nor g1080(n1138 ,n566 ,n756);
    nor g1081(n1137 ,n564 ,n754);
    nor g1082(n1136 ,n565 ,n766);
    nor g1083(n1135 ,n567 ,n750);
    nor g1084(n1134 ,n567 ,n754);
    nor g1085(n1133 ,n566 ,n754);
    nor g1086(n1132 ,n565 ,n754);
    nor g1087(n1131 ,n566 ,n750);
    nor g1088(n1130 ,n564 ,n758);
    nor g1089(n1129 ,n567 ,n758);
    nor g1090(n1128 ,n566 ,n758);
    nor g1091(n1127 ,n564 ,n780);
    nor g1092(n1126 ,n565 ,n758);
    nor g1093(n1125 ,n564 ,n760);
    nor g1094(n1124 ,n567 ,n780);
    nor g1095(n1123 ,n567 ,n760);
    nor g1096(n1122 ,n564 ,n762);
    nor g1097(n1121 ,n567 ,n762);
    nor g1098(n1120 ,n564 ,n756);
    nor g1099(n1119 ,n566 ,n760);
    nor g1100(n1118 ,n567 ,n756);
    nor g1101(n1117 ,n566 ,n762);
    nor g1102(n1116 ,n565 ,n756);
    nor g1103(n1115 ,n565 ,n762);
    nor g1104(n1114 ,n566 ,n780);
    nor g1105(n1113 ,n565 ,n760);
    nor g1106(n1112 ,n564 ,n764);
    nor g1107(n1111 ,n567 ,n764);
    nor g1108(n1110 ,n566 ,n764);
    nor g1109(n1109 ,n565 ,n780);
    nor g1110(n1108 ,n565 ,n764);
    nor g1111(n1107 ,n564 ,n770);
    nor g1112(n1106 ,n567 ,n770);
    nor g1113(n1105 ,n567 ,n778);
    nor g1114(n1104 ,n566 ,n778);
    nor g1115(n1103 ,n565 ,n778);
    nor g1116(n1102 ,n566 ,n770);
    nor g1117(n1101 ,n565 ,n770);
    nor g1118(n1100 ,n564 ,n774);
    nor g1119(n1099 ,n567 ,n774);
    nor g1120(n1098 ,n564 ,n772);
    nor g1121(n1097 ,n567 ,n772);
    nor g1122(n1096 ,n566 ,n774);
    nor g1123(n1095 ,n565 ,n774);
    nor g1124(n1094 ,n564 ,n768);
    nor g1125(n1093 ,n567 ,n768);
    nor g1126(n1092 ,n566 ,n772);
    nor g1127(n1091 ,n566 ,n768);
    nor g1128(n1090 ,n565 ,n768);
    nor g1129(n1089 ,n565 ,n750);
    nor g1130(n1088 ,n565 ,n772);
    nor g1131(n1087 ,n564 ,n750);
    nor g1132(n1086 ,n564 ,n752);
    nor g1133(n1085 ,n567 ,n752);
    nor g1134(n1084 ,n564 ,n778);
    nor g1135(n1083 ,n564 ,n766);
    nor g1136(n1082 ,n567 ,n766);
    nor g1137(n1081 ,n566 ,n752);
    nor g1138(n1080 ,n565 ,n752);
    or g1139(n1079 ,n956 ,n955);
    or g1140(n1078 ,n702 ,n747);
    or g1141(n1077 ,n715 ,n887);
    xor g1142(n1076 ,n26[0] ,n534);
    or g1143(n1075 ,n950 ,n798);
    or g1144(n1074 ,n682 ,n855);
    or g1145(n1073 ,n795 ,n945);
    or g1146(n1072 ,n809 ,n944);
    or g1147(n1071 ,n825 ,n822);
    or g1148(n1070 ,n908 ,n797);
    or g1149(n1069 ,n878 ,n927);
    or g1150(n1068 ,n900 ,n933);
    or g1151(n1067 ,n935 ,n790);
    or g1152(n1066 ,n876 ,n842);
    or g1153(n1065 ,n932 ,n942);
    or g1154(n1064 ,n720 ,n721);
    or g1155(n1063 ,n881 ,n865);
    or g1156(n1062 ,n854 ,n867);
    nor g1157(n1061 ,n784 ,n782);
    or g1158(n1060 ,n718 ,n922);
    or g1159(n1059 ,n905 ,n872);
    or g1160(n1058 ,n916 ,n729);
    or g1161(n1057 ,n717 ,n677);
    or g1162(n1056 ,n915 ,n835);
    or g1163(n1055 ,n909 ,n693);
    or g1164(n1054 ,n929 ,n725);
    or g1165(n1053 ,n681 ,n949);
    or g1166(n1052 ,n802 ,n726);
    or g1167(n1051 ,n918 ,n678);
    or g1168(n1050 ,n712 ,n896);
    or g1169(n1049 ,n938 ,n892);
    or g1170(n1048 ,n857 ,n799);
    or g1171(n1047 ,n953 ,n940);
    or g1172(n1046 ,n868 ,n858);
    or g1173(n1045 ,n706 ,n697);
    or g1174(n1044 ,n946 ,n948);
    or g1175(n1043 ,n947 ,n897);
    or g1176(n1042 ,n888 ,n815);
    or g1177(n1041 ,n704 ,n875);
    or g1178(n1040 ,n812 ,n882);
    or g1179(n1039 ,n931 ,n856);
    or g1180(n1038 ,n886 ,n869);
    or g1181(n1037 ,n690 ,n707);
    or g1182(n1036 ,n924 ,n814);
    or g1183(n1035 ,n831 ,n880);
    or g1184(n1034 ,n860 ,n864);
    or g1185(n1033 ,n852 ,n930);
    or g1186(n1032 ,n870 ,n851);
    or g1187(n1031 ,n846 ,n926);
    nor g1188(n1030 ,n1 ,n616);
    or g1189(n1029 ,n939 ,n827);
    or g1190(n1028 ,n843 ,n824);
    or g1191(n1027 ,n941 ,n819);
    or g1192(n1026 ,n688 ,n665);
    or g1193(n1025 ,n913 ,n917);
    or g1194(n1024 ,n834 ,n891);
    or g1195(n1023 ,n879 ,n885);
    or g1196(n1022 ,n808 ,n807);
    nor g1197(n1021 ,n1 ,n615);
    nor g1198(n1020 ,n1 ,n613);
    nor g1199(n1019 ,n1 ,n614);
    nor g1200(n1018 ,n1 ,n605);
    or g1201(n1017 ,n746 ,n849);
    nor g1202(n1016 ,n1 ,n601);
    nor g1203(n1015 ,n1 ,n617);
    or g1204(n1014 ,n687 ,n920);
    nor g1205(n1013 ,n1 ,n609);
    or g1206(n1012 ,n793 ,n832);
    or g1207(n1011 ,n664 ,n668);
    or g1208(n1010 ,n742 ,n666);
    or g1209(n1009 ,n740 ,n696);
    or g1210(n1008 ,n741 ,n739);
    or g1211(n1007 ,n889 ,n736);
    or g1212(n1006 ,n735 ,n734);
    or g1213(n1005 ,n733 ,n732);
    or g1214(n1004 ,n730 ,n743);
    or g1215(n1003 ,n728 ,n952);
    or g1216(n1002 ,n957 ,n727);
    or g1217(n1001 ,n691 ,n829);
    or g1218(n1000 ,n884 ,n679);
    or g1219(n999 ,n724 ,n806);
    or g1220(n998 ,n813 ,n723);
    or g1221(n997 ,n737 ,n811);
    or g1222(n996 ,n821 ,n719);
    or g1223(n995 ,n826 ,n823);
    or g1224(n994 ,n844 ,n839);
    or g1225(n993 ,n695 ,n792);
    or g1226(n992 ,n686 ,n838);
    or g1227(n991 ,n714 ,n791);
    or g1228(n990 ,n862 ,n796);
    or g1229(n989 ,n745 ,n841);
    or g1230(n988 ,n711 ,n866);
    or g1231(n987 ,n859 ,n850);
    or g1232(n986 ,n853 ,n709);
    or g1233(n985 ,n708 ,n861);
    or g1234(n984 ,n667 ,n951);
    or g1235(n983 ,n890 ,n919);
    or g1236(n982 ,n903 ,n901);
    or g1237(n981 ,n701 ,n912);
    or g1238(n980 ,n817 ,n700);
    or g1239(n979 ,n923 ,n902);
    or g1240(n978 ,n699 ,n863);
    or g1241(n977 ,n894 ,n898);
    or g1242(n976 ,n738 ,n836);
    or g1243(n975 ,n673 ,n694);
    or g1244(n974 ,n692 ,n883);
    or g1245(n973 ,n914 ,n899);
    or g1246(n972 ,n748 ,n710);
    or g1247(n971 ,n680 ,n685);
    or g1248(n970 ,n731 ,n937);
    or g1249(n969 ,n689 ,n936);
    or g1250(n968 ,n803 ,n800);
    or g1251(n967 ,n749 ,n789);
    or g1252(n966 ,n911 ,n934);
    or g1253(n965 ,n684 ,n818);
    or g1254(n964 ,n845 ,n910);
    or g1255(n963 ,n906 ,n830);
    or g1256(n962 ,n670 ,n804);
    or g1257(n961 ,n676 ,n874);
    or g1258(n960 ,n877 ,n928);
    or g1259(n959 ,n893 ,n895);
    or g1260(n958 ,n683 ,n671);
    nor g1261(n1208 ,n662 ,n602);
    nor g1262(n1207 ,n659 ,n599);
    nor g1263(n1206 ,n656 ,n603);
    nor g1264(n1205 ,n657 ,n612);
    nor g1265(n1204 ,n652 ,n620);
    nor g1266(n1203 ,n661 ,n611);
    nor g1267(n1202 ,n653 ,n608);
    nor g1268(n1201 ,n660 ,n607);
    nor g1269(n1200 ,n658 ,n604);
    nor g1270(n1199 ,n655 ,n610);
    nor g1271(n1198 ,n654 ,n619);
    nor g1272(n957 ,n386 ,n560);
    nor g1273(n956 ,n342 ,n589);
    nor g1274(n955 ,n433 ,n555);
    nor g1275(n954 ,n205 ,n558);
    nor g1276(n953 ,n227 ,n559);
    nor g1277(n952 ,n485 ,n586);
    nor g1278(n951 ,n375 ,n562);
    nor g1279(n950 ,n273 ,n588);
    nor g1280(n949 ,n188 ,n561);
    nor g1281(n948 ,n481 ,n555);
    nor g1282(n947 ,n251 ,n563);
    nor g1283(n946 ,n456 ,n589);
    nor g1284(n945 ,n234 ,n590);
    nor g1285(n944 ,n443 ,n555);
    nor g1286(n943 ,n463 ,n558);
    nor g1287(n942 ,n255 ,n555);
    nor g1288(n941 ,n427 ,n559);
    nor g1289(n940 ,n435 ,n562);
    nor g1290(n939 ,n453 ,n560);
    nor g1291(n938 ,n174 ,n559);
    nor g1292(n937 ,n396 ,n568);
    nor g1293(n936 ,n353 ,n568);
    nor g1294(n935 ,n192 ,n557);
    nor g1295(n934 ,n181 ,n555);
    nor g1296(n933 ,n442 ,n562);
    nor g1297(n932 ,n354 ,n589);
    nor g1298(n931 ,n418 ,n559);
    nor g1299(n930 ,n274 ,n586);
    nor g1300(n929 ,n490 ,n563);
    nor g1301(n928 ,n423 ,n586);
    nor g1302(n927 ,n399 ,n561);
    nor g1303(n926 ,n206 ,n590);
    nor g1304(n925 ,n250 ,n558);
    nor g1305(n924 ,n493 ,n557);
    nor g1306(n923 ,n259 ,n563);
    nor g1307(n922 ,n422 ,n555);
    nor g1308(n921 ,n380 ,n558);
    nor g1309(n920 ,n491 ,n587);
    nor g1310(n919 ,n374 ,n562);
    nor g1311(n918 ,n182 ,n559);
    nor g1312(n917 ,n476 ,n561);
    nor g1313(n916 ,n376 ,n560);
    nor g1314(n915 ,n248 ,n554);
    nor g1315(n914 ,n367 ,n554);
    nor g1316(n913 ,n432 ,n560);
    nor g1317(n912 ,n496 ,n562);
    nor g1318(n911 ,n403 ,n589);
    nor g1319(n910 ,n489 ,n586);
    nor g1320(n909 ,n439 ,n589);
    nor g1321(n908 ,n335 ,n559);
    nor g1322(n907 ,n238 ,n556);
    nor g1323(n906 ,n461 ,n560);
    nor g1324(n905 ,n401 ,n563);
    nor g1325(n904 ,n177 ,n558);
    nor g1326(n903 ,n180 ,n589);
    nor g1327(n902 ,n494 ,n586);
    nor g1328(n901 ,n245 ,n555);
    nor g1329(n900 ,n398 ,n559);
    nor g1330(n899 ,n253 ,n568);
    nor g1331(n898 ,n415 ,n587);
    nor g1332(n897 ,n373 ,n586);
    nor g1333(n896 ,n488 ,n587);
    nor g1334(n895 ,n408 ,n568);
    nor g1335(n894 ,n175 ,n557);
    nor g1336(n893 ,n328 ,n554);
    nor g1337(n892 ,n196 ,n562);
    nor g1338(n891 ,n469 ,n555);
    nor g1339(n890 ,n244 ,n559);
    nor g1340(n889 ,n212 ,n589);
    nor g1341(n888 ,n464 ,n560);
    nor g1342(n887 ,n497 ,n561);
    nor g1343(n886 ,n265 ,n554);
    nor g1344(n885 ,n249 ,n590);
    nor g1345(n884 ,n330 ,n557);
    nor g1346(n883 ,n260 ,n562);
    nor g1347(n882 ,n479 ,n590);
    nor g1348(n881 ,n269 ,n557);
    nor g1349(n880 ,n471 ,n590);
    nor g1350(n879 ,n387 ,n588);
    nor g1351(n878 ,n329 ,n560);
    nor g1352(n877 ,n345 ,n563);
    nor g1353(n876 ,n230 ,n588);
    nor g1354(n875 ,n458 ,n587);
    nor g1355(n874 ,n409 ,n555);
    nor g1356(n873 ,n189 ,n556);
    nor g1357(n872 ,n378 ,n586);
    nor g1358(n871 ,n220 ,n556);
    nor g1359(n870 ,n262 ,n554);
    nor g1360(n869 ,n199 ,n568);
    nor g1361(n868 ,n207 ,n589);
    nor g1362(n867 ,n420 ,n561);
    nor g1363(n866 ,n452 ,n562);
    nor g1364(n865 ,n242 ,n587);
    nor g1365(n864 ,n467 ,n590);
    nor g1366(n863 ,n500 ,n561);
    nor g1367(n862 ,n334 ,n563);
    nor g1368(n861 ,n462 ,n561);
    nor g1369(n860 ,n240 ,n588);
    nor g1370(n859 ,n176 ,n554);
    nor g1371(n858 ,n410 ,n555);
    nor g1372(n857 ,n449 ,n588);
    nor g1373(n856 ,n473 ,n562);
    nor g1374(n855 ,n209 ,n586);
    nor g1375(n854 ,n224 ,n560);
    nor g1376(n853 ,n271 ,n563);
    nor g1377(n852 ,n178 ,n563);
    nor g1378(n851 ,n336 ,n568);
    nor g1379(n850 ,n392 ,n568);
    nor g1380(n849 ,n268 ,n568);
    nor g1381(n848 ,n225 ,n558);
    nor g1382(n847 ,n419 ,n558);
    nor g1383(n846 ,n397 ,n588);
    nor g1384(n845 ,n213 ,n563);
    nor g1385(n844 ,n377 ,n560);
    nor g1386(n843 ,n276 ,n563);
    nor g1387(n842 ,n355 ,n590);
    nor g1388(n841 ,n237 ,n555);
    nor g1389(n840 ,n455 ,n558);
    nor g1390(n839 ,n272 ,n561);
    nor g1391(n838 ,n412 ,n587);
    nor g1392(n837 ,n215 ,n556);
    nor g1393(n836 ,n486 ,n586);
    nor g1394(n835 ,n444 ,n568);
    nor g1395(n834 ,n362 ,n589);
    nor g1396(n833 ,n350 ,n556);
    nor g1397(n832 ,n478 ,n590);
    nor g1398(n831 ,n228 ,n588);
    nor g1399(n830 ,n190 ,n561);
    nor g1400(n829 ,n333 ,n587);
    nor g1401(n828 ,n356 ,n556);
    nor g1402(n827 ,n231 ,n561);
    nor g1403(n826 ,n246 ,n563);
    nor g1404(n825 ,n413 ,n554);
    nor g1405(n824 ,n216 ,n586);
    nor g1406(n823 ,n402 ,n586);
    nor g1407(n822 ,n381 ,n568);
    nor g1408(n821 ,n424 ,n554);
    nor g1409(n820 ,n351 ,n558);
    nor g1410(n819 ,n487 ,n562);
    nor g1411(n818 ,n236 ,n562);
    nor g1412(n817 ,n451 ,n554);
    nor g1413(n816 ,n266 ,n558);
    nor g1414(n815 ,n352 ,n561);
    nor g1415(n814 ,n197 ,n587);
    nor g1416(n813 ,n232 ,n588);
    nor g1417(n812 ,n472 ,n588);
    nor g1418(n811 ,n277 ,n555);
    nor g1419(n810 ,n201 ,n556);
    nor g1420(n809 ,n390 ,n589);
    nor g1421(n808 ,n445 ,n557);
    nor g1422(n807 ,n384 ,n587);
    nor g1423(n806 ,n263 ,n587);
    nor g1424(n805 ,n414 ,n556);
    nor g1425(n804 ,n229 ,n590);
    nor g1426(n803 ,n267 ,n588);
    nor g1427(n802 ,n360 ,n554);
    nor g1428(n801 ,n448 ,n556);
    nor g1429(n800 ,n338 ,n590);
    nor g1430(n799 ,n388 ,n590);
    nor g1431(n798 ,n363 ,n590);
    nor g1432(n797 ,n256 ,n562);
    nor g1433(n796 ,n368 ,n586);
    nor g1434(n795 ,n219 ,n588);
    nor g1435(n794 ,n340 ,n556);
    nor g1436(n793 ,n436 ,n588);
    nor g1437(n792 ,n480 ,n587);
    nor g1438(n791 ,n191 ,n587);
    nor g1439(n790 ,n447 ,n587);
    nor g1440(n789 ,n411 ,n590);
    or g1441(n788 ,n152 ,n571);
    not g1442(n785 ,n784);
    not g1443(n783 ,n782);
    not g1444(n780 ,n781);
    not g1445(n778 ,n779);
    not g1446(n776 ,n777);
    not g1447(n774 ,n775);
    not g1448(n772 ,n773);
    not g1449(n770 ,n771);
    not g1450(n768 ,n769);
    not g1451(n766 ,n767);
    not g1452(n764 ,n765);
    not g1453(n762 ,n763);
    not g1454(n760 ,n761);
    not g1455(n758 ,n759);
    not g1456(n756 ,n757);
    not g1457(n754 ,n755);
    not g1458(n752 ,n753);
    not g1459(n750 ,n751);
    nor g1460(n749 ,n394 ,n588);
    nor g1461(n748 ,n247 ,n563);
    nor g1462(n747 ,n187 ,n568);
    nor g1463(n746 ,n339 ,n554);
    nor g1464(n745 ,n429 ,n589);
    nor g1465(n744 ,n371 ,n556);
    nor g1466(n743 ,n347 ,n568);
    nor g1467(n742 ,n404 ,n557);
    nor g1468(n741 ,n465 ,n588);
    nor g1469(n740 ,n477 ,n588);
    nor g1470(n739 ,n474 ,n590);
    nor g1471(n738 ,n440 ,n563);
    nor g1472(n737 ,n195 ,n589);
    nor g1473(n736 ,n400 ,n555);
    nor g1474(n735 ,n468 ,n557);
    nor g1475(n734 ,n341 ,n587);
    nor g1476(n733 ,n186 ,n559);
    nor g1477(n732 ,n454 ,n562);
    nor g1478(n731 ,n501 ,n554);
    nor g1479(n730 ,n194 ,n554);
    nor g1480(n729 ,n365 ,n561);
    nor g1481(n728 ,n475 ,n563);
    nor g1482(n727 ,n241 ,n561);
    nor g1483(n726 ,n372 ,n568);
    nor g1484(n725 ,n243 ,n586);
    nor g1485(n724 ,n343 ,n557);
    nor g1486(n723 ,n437 ,n590);
    nor g1487(n722 ,n222 ,n558);
    nor g1488(n721 ,n421 ,n562);
    nor g1489(n720 ,n382 ,n559);
    nor g1490(n719 ,n457 ,n568);
    nor g1491(n718 ,n450 ,n589);
    nor g1492(n717 ,n466 ,n559);
    nor g1493(n716 ,n239 ,n558);
    nor g1494(n715 ,n498 ,n560);
    nor g1495(n714 ,n332 ,n557);
    nor g1496(n713 ,n379 ,n558);
    nor g1497(n712 ,n235 ,n557);
    nor g1498(n711 ,n428 ,n559);
    nor g1499(n710 ,n434 ,n586);
    nor g1500(n709 ,n358 ,n586);
    nor g1501(n708 ,n483 ,n560);
    nor g1502(n707 ,n357 ,n586);
    nor g1503(n706 ,n492 ,n560);
    nor g1504(n705 ,n173 ,n556);
    nor g1505(n704 ,n369 ,n557);
    nor g1506(n703 ,n257 ,n558);
    nor g1507(n702 ,n417 ,n554);
    nor g1508(n701 ,n446 ,n559);
    nor g1509(n700 ,n221 ,n568);
    nor g1510(n699 ,n214 ,n560);
    nor g1511(n698 ,n385 ,n556);
    nor g1512(n697 ,n204 ,n561);
    nor g1513(n696 ,n208 ,n590);
    nor g1514(n695 ,n270 ,n557);
    nor g1515(n694 ,n430 ,n555);
    nor g1516(n693 ,n405 ,n555);
    nor g1517(n692 ,n364 ,n559);
    nor g1518(n691 ,n203 ,n557);
    nor g1519(n690 ,n226 ,n563);
    nor g1520(n689 ,n499 ,n554);
    nor g1521(n688 ,n264 ,n554);
    nor g1522(n687 ,n183 ,n557);
    nor g1523(n686 ,n502 ,n557);
    nor g1524(n685 ,n395 ,n561);
    nor g1525(n684 ,n211 ,n559);
    nor g1526(n683 ,n407 ,n560);
    nor g1527(n682 ,n391 ,n563);
    nor g1528(n681 ,n366 ,n560);
    nor g1529(n680 ,n441 ,n560);
    nor g1530(n679 ,n459 ,n587);
    nor g1531(n678 ,n223 ,n562);
    nor g1532(n677 ,n393 ,n562);
    nor g1533(n676 ,n348 ,n589);
    nor g1534(n675 ,n438 ,n558);
    nor g1535(n674 ,n349 ,n556);
    nor g1536(n673 ,n416 ,n589);
    nor g1537(n672 ,n406 ,n556);
    nor g1538(n671 ,n431 ,n561);
    nor g1539(n670 ,n200 ,n588);
    nor g1540(n669 ,n185 ,n558);
    nor g1541(n668 ,n359 ,n555);
    nor g1542(n667 ,n425 ,n559);
    nor g1543(n666 ,n331 ,n587);
    nor g1544(n665 ,n202 ,n568);
    nor g1545(n664 ,n184 ,n589);
    nor g1546(n663 ,n275 ,n556);
    nor g1547(n662 ,n158 ,n552);
    nor g1548(n661 ,n163 ,n552);
    nor g1549(n660 ,n166 ,n552);
    nor g1550(n659 ,n161 ,n552);
    nor g1551(n658 ,n157 ,n552);
    nor g1552(n657 ,n162 ,n552);
    nor g1553(n656 ,n170 ,n552);
    nor g1554(n655 ,n165 ,n552);
    nor g1555(n654 ,n164 ,n552);
    nor g1556(n653 ,n168 ,n552);
    nor g1557(n652 ,n159 ,n552);
    nor g1558(n651 ,n294 ,n550);
    nor g1559(n650 ,n310 ,n550);
    nor g1560(n649 ,n306 ,n550);
    nor g1561(n648 ,n308 ,n550);
    nor g1562(n647 ,n301 ,n550);
    nor g1563(n646 ,n303 ,n550);
    nor g1564(n645 ,n287 ,n550);
    nor g1565(n644 ,n309 ,n550);
    nor g1566(n643 ,n279 ,n550);
    nor g1567(n642 ,n288 ,n550);
    nor g1568(n641 ,n305 ,n550);
    nor g1569(n640 ,n281 ,n550);
    nor g1570(n639 ,n290 ,n550);
    nor g1571(n638 ,n304 ,n550);
    nor g1572(n637 ,n298 ,n550);
    nor g1573(n636 ,n210 ,n551);
    nor g1574(n635 ,n361 ,n551);
    nor g1575(n634 ,n389 ,n551);
    nor g1576(n633 ,n426 ,n551);
    nor g1577(n632 ,n179 ,n551);
    nor g1578(n631 ,n198 ,n551);
    nor g1579(n630 ,n344 ,n551);
    nor g1580(n629 ,n470 ,n551);
    nor g1581(n628 ,n484 ,n551);
    nor g1582(n627 ,n482 ,n551);
    nor g1583(n626 ,n252 ,n551);
    nor g1584(n625 ,n217 ,n551);
    nor g1585(n624 ,n370 ,n551);
    nor g1586(n623 ,n254 ,n551);
    nor g1587(n622 ,n218 ,n551);
    nor g1588(n621 ,n193 ,n551);
    nor g1589(n620 ,n544 ,n553);
    nor g1590(n619 ,n542 ,n553);
    or g1591(n618 ,n570 ,n598);
    nor g1592(n617 ,n585 ,n583);
    nor g1593(n616 ,n578 ,n536);
    nor g1594(n615 ,n574 ,n549);
    nor g1595(n614 ,n575 ,n580);
    nor g1596(n613 ,n572 ,n581);
    nor g1597(n612 ,n546 ,n553);
    nor g1598(n611 ,n548 ,n553);
    nor g1599(n610 ,n539 ,n553);
    nor g1600(n609 ,n577 ,n582);
    nor g1601(n608 ,n540 ,n553);
    nor g1602(n607 ,n547 ,n553);
    or g1603(n606 ,n598 ,n571);
    nor g1604(n605 ,n573 ,n579);
    nor g1605(n604 ,n541 ,n553);
    nor g1606(n603 ,n543 ,n553);
    nor g1607(n602 ,n545 ,n553);
    nor g1608(n601 ,n576 ,n584);
    or g1609(n600 ,n26[0] ,n570);
    nor g1610(n599 ,n538 ,n553);
    or g1611(n787 ,n1 ,n535);
    or g1612(n786 ,n1 ,n537);
    nor g1613(n784 ,n550 ,n553);
    nor g1614(n782 ,n550 ,n552);
    nor g1615(n781 ,n594 ,n593);
    nor g1616(n779 ,n596 ,n569);
    nor g1617(n777 ,n595 ,n592);
    nor g1618(n775 ,n594 ,n592);
    nor g1619(n773 ,n597 ,n569);
    nor g1620(n771 ,n594 ,n569);
    nor g1621(n769 ,n595 ,n593);
    nor g1622(n767 ,n596 ,n593);
    nor g1623(n765 ,n595 ,n569);
    nor g1624(n763 ,n597 ,n591);
    nor g1625(n761 ,n597 ,n593);
    nor g1626(n759 ,n595 ,n591);
    nor g1627(n757 ,n596 ,n591);
    nor g1628(n755 ,n596 ,n592);
    nor g1629(n753 ,n597 ,n592);
    nor g1630(n751 ,n594 ,n591);
    nor g1631(n585 ,n383 ,n529);
    nor g1632(n584 ,n300 ,n528);
    nor g1633(n583 ,n285 ,n528);
    nor g1634(n582 ,n291 ,n528);
    nor g1635(n581 ,n295 ,n526);
    nor g1636(n580 ,n293 ,n526);
    nor g1637(n579 ,n278 ,n526);
    nor g1638(n578 ,n337 ,n529);
    nor g1639(n577 ,n460 ,n529);
    nor g1640(n576 ,n346 ,n529);
    nor g1641(n575 ,n495 ,n527);
    nor g1642(n574 ,n233 ,n527);
    nor g1643(n573 ,n261 ,n527);
    nor g1644(n572 ,n258 ,n527);
    or g1645(n598 ,n509 ,n511);
    or g1646(n597 ,n141 ,n510);
    or g1647(n596 ,n141 ,n517);
    or g1648(n595 ,n141 ,n516);
    or g1649(n594 ,n141 ,n507);
    or g1650(n593 ,n133 ,n132);
    or g1651(n592 ,n131 ,n132);
    or g1652(n591 ,n130 ,n133);
    or g1653(n590 ,n512 ,n514);
    or g1654(n589 ,n531 ,n532);
    or g1655(n588 ,n532 ,n512);
    or g1656(n587 ,n532 ,n515);
    or g1657(n586 ,n515 ,n514);
    not g1658(n552 ,n553);
    not g1659(n550 ,n551);
    nor g1660(n549 ,n27[0] ,n526);
    xnor g1661(n548 ,n4[9] ,n29[9]);
    xnor g1662(n547 ,n4[13] ,n29[13]);
    xnor g1663(n546 ,n4[4] ,n29[4]);
    xnor g1664(n545 ,n4[6] ,n29[6]);
    xnor g1665(n544 ,n4[10] ,n29[10]);
    xnor g1666(n543 ,n4[7] ,n29[7]);
    xnor g1667(n542 ,n4[12] ,n29[12]);
    xnor g1668(n541 ,n4[14] ,n29[14]);
    xnor g1669(n540 ,n4[5] ,n29[5]);
    xnor g1670(n539 ,n4[11] ,n29[11]);
    xnor g1671(n538 ,n4[8] ,n29[8]);
    or g1672(n537 ,n527 ,n529);
    nor g1673(n536 ,n28[0] ,n528);
    or g1674(n535 ,n527 ,n528);
    nor g1675(n534 ,n527 ,n529);
    or g1676(n571 ,n503 ,n504);
    or g1677(n570 ,n26[5] ,n508);
    or g1678(n569 ,n131 ,n130);
    or g1679(n568 ,n531 ,n514);
    xnor g1680(n567 ,n4[1] ,n29[1]);
    xnor g1681(n566 ,n4[2] ,n29[2]);
    xnor g1682(n565 ,n4[3] ,n29[3]);
    xnor g1683(n564 ,n4[0] ,n29[0]);
    or g1684(n563 ,n530 ,n513);
    or g1685(n562 ,n533 ,n512);
    or g1686(n561 ,n530 ,n514);
    or g1687(n560 ,n513 ,n512);
    or g1688(n559 ,n531 ,n513);
    or g1689(n558 ,n531 ,n533);
    or g1690(n557 ,n533 ,n530);
    or g1691(n556 ,n532 ,n530);
    or g1692(n555 ,n533 ,n515);
    or g1693(n554 ,n515 ,n513);
    nor g1694(n553 ,n505 ,n506);
    nor g1695(n551 ,n1 ,n526);
    not g1696(n528 ,n529);
    not g1697(n526 ,n527);
    nor g1698(n525 ,n337 ,n1);
    nor g1699(n524 ,n383 ,n1);
    nor g1700(n523 ,n495 ,n1);
    nor g1701(n522 ,n346 ,n1);
    nor g1702(n521 ,n261 ,n1);
    nor g1703(n520 ,n258 ,n1);
    nor g1704(n519 ,n233 ,n1);
    nor g1705(n518 ,n460 ,n1);
    or g1706(n517 ,n315 ,n142);
    or g1707(n516 ,n142 ,n28[0]);
    or g1708(n533 ,n316 ,n144);
    or g1709(n532 ,n144 ,n27[0]);
    or g1710(n531 ,n143 ,n140);
    or g1711(n530 ,n143 ,n27[2]);
    nor g1712(n529 ,n141 ,n7);
    nor g1713(n527 ,n311 ,n6);
    or g1714(n511 ,n26[10] ,n26[11]);
    or g1715(n510 ,n315 ,n28[3]);
    or g1716(n509 ,n26[8] ,n26[9]);
    or g1717(n508 ,n26[6] ,n26[7]);
    or g1718(n507 ,n28[0] ,n28[3]);
    or g1719(n506 ,n29[1] ,n29[0]);
    or g1720(n505 ,n29[3] ,n29[2]);
    or g1721(n504 ,n26[14] ,n26[15]);
    or g1722(n503 ,n26[12] ,n26[13]);
    or g1723(n515 ,n140 ,n27[1]);
    or g1724(n514 ,n27[0] ,n27[3]);
    or g1725(n513 ,n316 ,n27[3]);
    or g1726(n512 ,n27[1] ,n27[2]);
    not g1727(n495 ,n24[2]);
    not g1728(n484 ,n5[6]);
    not g1729(n482 ,n5[14]);
    not g1730(n470 ,n5[7]);
    not g1731(n460 ,n25[3]);
    not g1732(n426 ,n5[10]);
    not g1733(n389 ,n5[15]);
    not g1734(n383 ,n25[2]);
    not g1735(n370 ,n5[12]);
    not g1736(n361 ,n5[5]);
    not g1737(n346 ,n25[1]);
    not g1738(n344 ,n5[8]);
    not g1739(n337 ,n25[0]);
    not g1740(n327 ,n26[5]);
    not g1741(n326 ,n26[8]);
    not g1742(n325 ,n26[11]);
    not g1743(n324 ,n26[6]);
    not g1744(n323 ,n26[13]);
    not g1745(n322 ,n26[14]);
    not g1746(n321 ,n26[1]);
    not g1747(n320 ,n26[2]);
    not g1748(n319 ,n26[3]);
    not g1749(n318 ,n28[1]);
    not g1750(n317 ,n28[2]);
    not g1751(n316 ,n27[0]);
    not g1752(n315 ,n28[0]);
    not g1753(n314 ,n2209);
    not g1754(n313 ,n2205);
    not g1755(n312 ,n2202);
    not g1756(n311 ,n3);
    not g1757(n310 ,n2185);
    not g1758(n309 ,n2192);
    not g1759(n308 ,n2194);
    not g1760(n307 ,n2206);
    not g1761(n306 ,n2183);
    not g1762(n305 ,n2191);
    not g1763(n304 ,n2188);
    not g1764(n303 ,n2180);
    not g1765(n302 ,n2199);
    not g1766(n301 ,n2181);
    not g1767(n300 ,n2212);
    not g1768(n299 ,n2208);
    not g1769(n298 ,n2187);
    not g1770(n297 ,n2198);
    not g1771(n296 ,n2201);
    not g1772(n295 ,n2215);
    not g1773(n294 ,n2184);
    not g1774(n293 ,n2214);
    not g1775(n292 ,n2195);
    not g1776(n291 ,n2210);
    not g1777(n290 ,n2189);
    not g1778(n289 ,n2207);
    not g1779(n288 ,n2182);
    not g1780(n287 ,n2186);
    not g1781(n286 ,n2196);
    not g1782(n285 ,n2211);
    not g1783(n284 ,n2204);
    not g1784(n283 ,n2197);
    not g1785(n282 ,n2203);
    not g1786(n281 ,n2193);
    not g1787(n280 ,n2200);
    not g1788(n279 ,n2190);
    not g1789(n278 ,n2213);
    not g1790(n261 ,n24[3]);
    not g1791(n258 ,n24[1]);
    not g1792(n254 ,n5[2]);
    not g1793(n252 ,n5[0]);
    not g1794(n233 ,n24[0]);
    not g1795(n218 ,n5[1]);
    not g1796(n217 ,n5[11]);
    not g1797(n210 ,n5[3]);
    not g1798(n198 ,n5[9]);
    not g1799(n193 ,n5[4]);
    not g1800(n179 ,n5[13]);
    not g1801(n172 ,n26[9]);
    not g1802(n171 ,n26[10]);
    not g1803(n170 ,n4[7]);
    not g1804(n169 ,n26[7]);
    not g1805(n168 ,n4[5]);
    not g1806(n167 ,n26[12]);
    not g1807(n166 ,n4[13]);
    not g1808(n165 ,n4[11]);
    not g1809(n164 ,n4[12]);
    not g1810(n163 ,n4[9]);
    not g1811(n162 ,n4[4]);
    not g1812(n161 ,n4[8]);
    not g1813(n160 ,n26[15]);
    not g1814(n159 ,n4[10]);
    not g1815(n158 ,n4[6]);
    not g1816(n157 ,n4[14]);
    not g1817(n156 ,n29[13]);
    not g1818(n155 ,n29[6]);
    not g1819(n154 ,n29[7]);
    not g1820(n153 ,n29[9]);
    not g1821(n152 ,n26[4]);
    not g1822(n151 ,n29[10]);
    not g1823(n150 ,n29[14]);
    not g1824(n149 ,n29[5]);
    not g1825(n148 ,n29[4]);
    not g1826(n147 ,n29[11]);
    not g1827(n146 ,n29[12]);
    not g1828(n145 ,n29[8]);
    not g1829(n144 ,n27[3]);
    not g1830(n143 ,n27[1]);
    not g1831(n142 ,n28[3]);
    not g1832(n141 ,n2);
    not g1833(n140 ,n27[2]);
    not g1834(n139 ,n29[1]);
    not g1835(n138 ,n29[2]);
    not g1836(n137 ,n29[3]);
    not g1837(n136 ,n29[0]);
    not g1838(n135 ,n4[15]);
    or g1839(n134 ,n26[1] ,n26[2]);
    or g1840(n133 ,n7 ,n28[1]);
    or g1841(n132 ,n28[2] ,n1);
    or g1842(n131 ,n318 ,n7);
    or g1843(n130 ,n317 ,n1);
    xor g1844(n2194 ,n26[15] ,n57);
    xor g1845(n2193 ,n26[14] ,n55);
    nor g1846(n57 ,n26[14] ,n56);
    xor g1847(n2192 ,n26[13] ,n53);
    not g1848(n56 ,n55);
    nor g1849(n55 ,n26[13] ,n54);
    xor g1850(n2191 ,n26[12] ,n51);
    not g1851(n54 ,n53);
    nor g1852(n53 ,n26[12] ,n52);
    xor g1853(n2190 ,n26[11] ,n49);
    not g1854(n52 ,n51);
    nor g1855(n51 ,n26[11] ,n50);
    xor g1856(n2189 ,n26[10] ,n47);
    not g1857(n50 ,n49);
    nor g1858(n49 ,n26[10] ,n48);
    xor g1859(n2188 ,n26[9] ,n45);
    not g1860(n48 ,n47);
    nor g1861(n47 ,n26[9] ,n46);
    xor g1862(n2187 ,n26[8] ,n43);
    not g1863(n46 ,n45);
    nor g1864(n45 ,n26[8] ,n44);
    xor g1865(n2186 ,n26[7] ,n41);
    not g1866(n44 ,n43);
    nor g1867(n43 ,n26[7] ,n42);
    xor g1868(n2185 ,n26[6] ,n39);
    not g1869(n42 ,n41);
    nor g1870(n41 ,n26[6] ,n40);
    xor g1871(n2184 ,n26[5] ,n37);
    not g1872(n40 ,n39);
    nor g1873(n39 ,n26[5] ,n38);
    xor g1874(n2183 ,n26[4] ,n35);
    not g1875(n38 ,n37);
    nor g1876(n37 ,n26[4] ,n36);
    xor g1877(n2182 ,n26[3] ,n33);
    not g1878(n36 ,n35);
    nor g1879(n35 ,n26[3] ,n34);
    xor g1880(n2181 ,n26[2] ,n31);
    not g1881(n34 ,n33);
    nor g1882(n33 ,n26[2] ,n32);
    xnor g1883(n2180 ,n26[1] ,n26[0]);
    not g1884(n32 ,n31);
    nor g1885(n31 ,n26[1] ,n26[0]);
    xor g1886(n2210 ,n28[3] ,n65);
    nor g1887(n2211 ,n64 ,n65);
    nor g1888(n65 ,n60 ,n63);
    nor g1889(n64 ,n28[2] ,n62);
    nor g1890(n2212 ,n62 ,n61);
    not g1891(n63 ,n62);
    nor g1892(n62 ,n58 ,n59);
    nor g1893(n61 ,n28[1] ,n28[0]);
    not g1894(n60 ,n28[2]);
    not g1895(n59 ,n28[0]);
    not g1896(n58 ,n28[1]);
    xor g1897(n2209 ,n26[15] ,n121);
    nor g1898(n2208 ,n120 ,n121);
    nor g1899(n121 ,n77 ,n119);
    nor g1900(n120 ,n26[14] ,n118);
    nor g1901(n2207 ,n117 ,n118);
    not g1902(n119 ,n118);
    nor g1903(n118 ,n67 ,n116);
    nor g1904(n117 ,n26[13] ,n115);
    nor g1905(n2206 ,n114 ,n115);
    not g1906(n116 ,n115);
    nor g1907(n115 ,n80 ,n113);
    nor g1908(n114 ,n26[12] ,n112);
    nor g1909(n2205 ,n111 ,n112);
    not g1910(n113 ,n112);
    nor g1911(n112 ,n76 ,n110);
    nor g1912(n111 ,n26[11] ,n109);
    nor g1913(n2204 ,n108 ,n109);
    not g1914(n110 ,n109);
    nor g1915(n109 ,n78 ,n107);
    nor g1916(n108 ,n26[10] ,n106);
    nor g1917(n2203 ,n105 ,n106);
    not g1918(n107 ,n106);
    nor g1919(n106 ,n75 ,n104);
    nor g1920(n105 ,n26[9] ,n103);
    nor g1921(n2202 ,n102 ,n103);
    not g1922(n104 ,n103);
    nor g1923(n103 ,n72 ,n101);
    nor g1924(n102 ,n26[8] ,n100);
    nor g1925(n2201 ,n99 ,n100);
    not g1926(n101 ,n100);
    nor g1927(n100 ,n73 ,n98);
    nor g1928(n99 ,n26[7] ,n97);
    nor g1929(n2200 ,n96 ,n97);
    not g1930(n98 ,n97);
    nor g1931(n97 ,n66 ,n95);
    nor g1932(n96 ,n26[6] ,n94);
    nor g1933(n2199 ,n93 ,n94);
    not g1934(n95 ,n94);
    nor g1935(n94 ,n71 ,n92);
    nor g1936(n93 ,n26[5] ,n91);
    nor g1937(n2198 ,n90 ,n91);
    not g1938(n92 ,n91);
    nor g1939(n91 ,n69 ,n89);
    nor g1940(n90 ,n26[4] ,n88);
    nor g1941(n2197 ,n87 ,n88);
    not g1942(n89 ,n88);
    nor g1943(n88 ,n68 ,n86);
    nor g1944(n87 ,n26[3] ,n85);
    nor g1945(n2196 ,n84 ,n85);
    not g1946(n86 ,n85);
    nor g1947(n85 ,n70 ,n83);
    nor g1948(n84 ,n26[2] ,n82);
    nor g1949(n2195 ,n82 ,n81);
    not g1950(n83 ,n82);
    nor g1951(n82 ,n74 ,n79);
    nor g1952(n81 ,n26[1] ,n26[0]);
    not g1953(n80 ,n26[12]);
    not g1954(n79 ,n26[0]);
    not g1955(n78 ,n26[10]);
    not g1956(n77 ,n26[14]);
    not g1957(n76 ,n26[11]);
    not g1958(n75 ,n26[9]);
    not g1959(n74 ,n26[1]);
    not g1960(n73 ,n26[7]);
    not g1961(n72 ,n26[8]);
    not g1962(n71 ,n26[5]);
    not g1963(n70 ,n26[2]);
    not g1964(n69 ,n26[4]);
    not g1965(n68 ,n26[3]);
    not g1966(n67 ,n26[13]);
    not g1967(n66 ,n26[6]);
    xor g1968(n2213 ,n27[3] ,n129);
    nor g1969(n2214 ,n128 ,n129);
    nor g1970(n129 ,n124 ,n127);
    nor g1971(n128 ,n27[2] ,n126);
    nor g1972(n2215 ,n126 ,n125);
    not g1973(n127 ,n126);
    nor g1974(n126 ,n122 ,n123);
    nor g1975(n125 ,n27[1] ,n27[0]);
    not g1976(n124 ,n27[2]);
    not g1977(n123 ,n27[0]);
    not g1978(n122 ,n27[1]);
    xor g1979(n3646 ,n28[1] ,n27[1]);
    or g1980(n29[3] ,n3617 ,n3636);
    or g1981(n29[7] ,n3614 ,n3628);
    or g1982(n29[9] ,n3609 ,n3629);
    or g1983(n29[2] ,n3615 ,n3635);
    or g1984(n29[1] ,n3612 ,n3633);
    or g1985(n29[8] ,n3603 ,n3637);
    or g1986(n29[0] ,n3611 ,n3631);
    or g1987(n29[6] ,n3610 ,n3632);
    or g1988(n29[5] ,n3607 ,n3630);
    or g1989(n29[4] ,n3605 ,n3634);
    or g1990(n29[11] ,n3608 ,n3604);
    or g1991(n29[10] ,n3616 ,n3613);
    or g1992(n29[12] ,n3569 ,n3606);
    or g1993(n3637 ,n3602 ,n3627);
    or g1994(n3636 ,n3590 ,n3626);
    or g1995(n3635 ,n3588 ,n3625);
    or g1996(n3634 ,n3579 ,n3618);
    or g1997(n3633 ,n3597 ,n3624);
    or g1998(n3632 ,n3582 ,n3621);
    or g1999(n3631 ,n3580 ,n3622);
    or g2000(n3630 ,n3581 ,n3619);
    or g2001(n3629 ,n3568 ,n3620);
    or g2002(n3628 ,n3571 ,n3623);
    nor g2003(n3627 ,n3541 ,n3559);
    nor g2004(n3626 ,n3546 ,n3551);
    nor g2005(n3625 ,n3544 ,n3558);
    nor g2006(n3624 ,n3547 ,n3557);
    nor g2007(n3623 ,n3542 ,n3556);
    nor g2008(n3622 ,n3543 ,n3555);
    nor g2009(n3621 ,n3540 ,n3554);
    nor g2010(n3620 ,n3538 ,n3552);
    nor g2011(n3619 ,n3539 ,n3553);
    nor g2012(n3618 ,n3545 ,n3550);
    or g2013(n3617 ,n3601 ,n3576);
    or g2014(n3616 ,n3563 ,n3598);
    or g2015(n3615 ,n3600 ,n3574);
    or g2016(n3614 ,n3589 ,n3599);
    or g2017(n3613 ,n3586 ,n3572);
    or g2018(n3612 ,n3587 ,n3573);
    or g2019(n3611 ,n3596 ,n3577);
    or g2020(n3610 ,n3595 ,n3570);
    or g2021(n3609 ,n3583 ,n3593);
    or g2022(n3608 ,n3584 ,n3594);
    or g2023(n3607 ,n3592 ,n3567);
    or g2024(n29[13] ,n3560 ,n3575);
    or g2025(n3606 ,n3562 ,n3585);
    or g2026(n3605 ,n3591 ,n3566);
    or g2027(n3604 ,n3561 ,n3565);
    or g2028(n3603 ,n3578 ,n3564);
    nor g2029(n3602 ,n3472 ,n3537);
    nor g2030(n3601 ,n3475 ,n3537);
    nor g2031(n3600 ,n3499 ,n3537);
    nor g2032(n3599 ,n3474 ,n3537);
    nor g2033(n3598 ,n3473 ,n3537);
    nor g2034(n3597 ,n3497 ,n3537);
    nor g2035(n3596 ,n3495 ,n3537);
    nor g2036(n3595 ,n3503 ,n3537);
    nor g2037(n3594 ,n3502 ,n3537);
    nor g2038(n3593 ,n3500 ,n3537);
    nor g2039(n3592 ,n3498 ,n3537);
    nor g2040(n3591 ,n3501 ,n3537);
    nor g2041(n3590 ,n3513 ,n3549);
    nor g2042(n3589 ,n3508 ,n3549);
    nor g2043(n3588 ,n3486 ,n3549);
    nor g2044(n3587 ,n3518 ,n3549);
    nor g2045(n3586 ,n3520 ,n3549);
    nor g2046(n3585 ,n3483 ,n3549);
    nor g2047(n3584 ,n3511 ,n3549);
    nor g2048(n3583 ,n3522 ,n3549);
    nor g2049(n3582 ,n3524 ,n3549);
    nor g2050(n3581 ,n3525 ,n3549);
    nor g2051(n3580 ,n3487 ,n3549);
    nor g2052(n3579 ,n3485 ,n3549);
    nor g2053(n3578 ,n3509 ,n3549);
    nor g2054(n3577 ,n3516 ,n3536);
    nor g2055(n3576 ,n3521 ,n3536);
    nor g2056(n3575 ,n3496 ,n3536);
    nor g2057(n3574 ,n3488 ,n3536);
    nor g2058(n3573 ,n3482 ,n3536);
    nor g2059(n3572 ,n3493 ,n3536);
    nor g2060(n3571 ,n3484 ,n3536);
    nor g2061(n3570 ,n3489 ,n3536);
    nor g2062(n3569 ,n3519 ,n3536);
    nor g2063(n3568 ,n3491 ,n3536);
    nor g2064(n3567 ,n3490 ,n3536);
    nor g2065(n3566 ,n3492 ,n3536);
    nor g2066(n3565 ,n3514 ,n3536);
    nor g2067(n3564 ,n3494 ,n3536);
    nor g2068(n3563 ,n3515 ,n3548);
    nor g2069(n3562 ,n3523 ,n3548);
    nor g2070(n29[14] ,n3512 ,n3548);
    nor g2071(n3561 ,n3517 ,n3548);
    nor g2072(n3560 ,n3510 ,n3548);
    or g2073(n3559 ,n3548 ,n3528);
    or g2074(n3558 ,n3548 ,n3535);
    or g2075(n3557 ,n3548 ,n3531);
    or g2076(n3556 ,n3548 ,n3534);
    or g2077(n3555 ,n3548 ,n3533);
    or g2078(n3554 ,n3548 ,n3530);
    or g2079(n3553 ,n3548 ,n3526);
    or g2080(n3552 ,n3548 ,n3532);
    or g2081(n3551 ,n3548 ,n3529);
    or g2082(n3550 ,n3548 ,n3527);
    nor g2083(n3547 ,n3477 ,n3475);
    nor g2084(n3546 ,n3476 ,n3498);
    nor g2085(n3545 ,n3480 ,n3503);
    nor g2086(n3544 ,n3504 ,n3501);
    nor g2087(n3543 ,n3506 ,n3499);
    nor g2088(n3542 ,n3479 ,n3500);
    nor g2089(n3541 ,n3507 ,n3473);
    nor g2090(n3540 ,n3505 ,n3472);
    nor g2091(n3539 ,n3481 ,n3474);
    nor g2092(n3538 ,n3478 ,n3502);
    or g2093(n3549 ,n3470 ,n2);
    or g2094(n3548 ,n3471 ,n3470);
    nor g2095(n3535 ,n3692 ,n30[4]);
    nor g2096(n3534 ,n3687 ,n30[9]);
    nor g2097(n3533 ,n3694 ,n30[2]);
    nor g2098(n3532 ,n3685 ,n30[11]);
    nor g2099(n3531 ,n3693 ,n30[3]);
    nor g2100(n3530 ,n3688 ,n30[8]);
    nor g2101(n3529 ,n3691 ,n30[5]);
    nor g2102(n3528 ,n3686 ,n30[10]);
    nor g2103(n3527 ,n3690 ,n30[6]);
    nor g2104(n3526 ,n3689 ,n30[7]);
    or g2105(n3537 ,n3471 ,n3);
    or g2106(n3536 ,n2 ,n3);
    not g2107(n3525 ,n3654);
    not g2108(n3524 ,n3655);
    not g2109(n3523 ,n3642);
    not g2110(n3522 ,n3658);
    not g2111(n3521 ,n3665);
    not g2112(n3520 ,n3659);
    not g2113(n3519 ,n3674);
    not g2114(n3518 ,n3650);
    not g2115(n3517 ,n3641);
    not g2116(n3516 ,n3662);
    not g2117(n3515 ,n3640);
    not g2118(n3514 ,n3673);
    not g2119(n3513 ,n3652);
    not g2120(n3512 ,n3644);
    not g2121(n3511 ,n3660);
    not g2122(n3510 ,n3643);
    not g2123(n3509 ,n3657);
    not g2124(n3508 ,n3656);
    not g2125(n3507 ,n3686);
    not g2126(n3506 ,n3694);
    not g2127(n3505 ,n3688);
    not g2128(n3504 ,n3692);
    not g2129(n3503 ,n30[6]);
    not g2130(n3502 ,n30[11]);
    not g2131(n3501 ,n30[4]);
    not g2132(n3500 ,n30[9]);
    not g2133(n3499 ,n30[2]);
    not g2134(n3498 ,n30[5]);
    not g2135(n3497 ,n3639);
    not g2136(n3496 ,n3675);
    not g2137(n3495 ,n3638);
    not g2138(n3494 ,n3670);
    not g2139(n3493 ,n3672);
    not g2140(n3492 ,n3666);
    not g2141(n3491 ,n3671);
    not g2142(n3490 ,n3667);
    not g2143(n3489 ,n3668);
    not g2144(n3488 ,n3664);
    not g2145(n3487 ,n3649);
    not g2146(n3486 ,n3651);
    not g2147(n3485 ,n3653);
    not g2148(n3484 ,n3669);
    not g2149(n3483 ,n3661);
    not g2150(n3482 ,n3663);
    not g2151(n3481 ,n3689);
    not g2152(n3480 ,n3690);
    not g2153(n3479 ,n3687);
    not g2154(n3478 ,n3685);
    not g2155(n3477 ,n3693);
    not g2156(n3476 ,n3691);
    not g2157(n3475 ,n30[3]);
    not g2158(n3474 ,n30[7]);
    not g2159(n3473 ,n30[10]);
    not g2160(n3472 ,n30[8]);
    not g2161(n3471 ,n2);
    not g2162(n3470 ,n3);
    xor g2163(n3645 ,n28[0] ,n27[0]);
    xor g2164(n3647 ,n28[2] ,n27[2]);
    xor g2165(n3648 ,n28[3] ,n27[3]);
    or g2166(n3675 ,n2469 ,n2564);
    xnor g2167(n3674 ,n2480 ,n2563);
    nor g2168(n2564 ,n2473 ,n2563);
    nor g2169(n2563 ,n2504 ,n2562);
    xor g2170(n3673 ,n2513 ,n2561);
    nor g2171(n2562 ,n2503 ,n2561);
    nor g2172(n2561 ,n2524 ,n2560);
    xnor g2173(n3672 ,n2529 ,n2559);
    nor g2174(n2560 ,n2523 ,n2559);
    nor g2175(n2559 ,n2547 ,n2558);
    xnor g2176(n3671 ,n2549 ,n2557);
    nor g2177(n2558 ,n2548 ,n2557);
    nor g2178(n2557 ,n2536 ,n2556);
    xor g2179(n3670 ,n2545 ,n2555);
    nor g2180(n2556 ,n2539 ,n2555);
    nor g2181(n2555 ,n2533 ,n2554);
    xor g2182(n3669 ,n2544 ,n2553);
    nor g2183(n2554 ,n2538 ,n2553);
    nor g2184(n2553 ,n2532 ,n2552);
    xor g2185(n3668 ,n2543 ,n2551);
    nor g2186(n2552 ,n2541 ,n2551);
    nor g2187(n2551 ,n2537 ,n2550);
    xor g2188(n3667 ,n2542 ,n2546);
    nor g2189(n2550 ,n2540 ,n2546);
    xnor g2190(n2549 ,n2534 ,n2495);
    xnor g2191(n3666 ,n2530 ,n2522);
    nor g2192(n2548 ,n2496 ,n2534);
    nor g2193(n2547 ,n2495 ,n2535);
    nor g2194(n2546 ,n2525 ,n2531);
    xnor g2195(n2545 ,n2516 ,n2527);
    xnor g2196(n2544 ,n2518 ,n2509);
    xnor g2197(n2543 ,n2520 ,n2499);
    xnor g2198(n2542 ,n2514 ,n2511);
    nor g2199(n2541 ,n2500 ,n2521);
    nor g2200(n2540 ,n2512 ,n2515);
    nor g2201(n2539 ,n2528 ,n2517);
    nor g2202(n2538 ,n2510 ,n2519);
    nor g2203(n2537 ,n2511 ,n2514);
    nor g2204(n2536 ,n2527 ,n2516);
    not g2205(n2535 ,n2534);
    xor g2206(n3665 ,n2494 ,n2492);
    nor g2207(n2533 ,n2509 ,n2518);
    nor g2208(n2532 ,n2499 ,n2520);
    nor g2209(n2531 ,n2526 ,n2522);
    xnor g2210(n2530 ,n2501 ,n2474);
    xnor g2211(n2529 ,n2497 ,n2507);
    xnor g2212(n2534 ,n2493 ,n2433);
    not g2213(n2528 ,n2527);
    nor g2214(n2526 ,n2475 ,n2501);
    nor g2215(n2525 ,n2474 ,n2502);
    nor g2216(n2524 ,n2507 ,n2498);
    nor g2217(n2523 ,n2508 ,n2497);
    nor g2218(n2527 ,n2486 ,n2506);
    not g2219(n2521 ,n2520);
    not g2220(n2519 ,n2518);
    not g2221(n2517 ,n2516);
    not g2222(n2515 ,n2514);
    xnor g2223(n2513 ,n2454 ,n2483);
    nor g2224(n2522 ,n2487 ,n2505);
    xnor g2225(n2520 ,n2478 ,n2460);
    xnor g2226(n2518 ,n2476 ,n2452);
    xnor g2227(n2516 ,n2477 ,n2463);
    xnor g2228(n2514 ,n2479 ,n2458);
    not g2229(n2512 ,n2511);
    not g2230(n2510 ,n2509);
    not g2231(n2508 ,n2507);
    nor g2232(n2506 ,n2439 ,n2490);
    nor g2233(n2505 ,n2492 ,n2485);
    nor g2234(n2504 ,n2454 ,n2483);
    nor g2235(n2503 ,n2455 ,n2484);
    nor g2236(n2511 ,n2429 ,n2491);
    nor g2237(n2509 ,n2464 ,n2482);
    nor g2238(n2507 ,n2466 ,n2489);
    not g2239(n2502 ,n2501);
    not g2240(n2500 ,n2499);
    not g2241(n2498 ,n2497);
    not g2242(n2496 ,n2495);
    xor g2243(n3664 ,n2448 ,n2391);
    xnor g2244(n2494 ,n2456 ,n2405);
    xnor g2245(n2493 ,n2461 ,n2367);
    xnor g2246(n2501 ,n2430 ,n2459);
    nor g2247(n2499 ,n2450 ,n2481);
    xnor g2248(n2497 ,n2449 ,n2440);
    nor g2249(n2495 ,n2451 ,n2488);
    nor g2250(n2491 ,n2428 ,n2459);
    nor g2251(n2490 ,n2344 ,n2453);
    nor g2252(n2489 ,n2471 ,n2462);
    nor g2253(n2488 ,n2468 ,n2463);
    nor g2254(n2487 ,n2406 ,n2457);
    nor g2255(n2486 ,n2343 ,n2452);
    nor g2256(n2485 ,n2405 ,n2456);
    nor g2257(n2492 ,n2443 ,n2467);
    not g2258(n2484 ,n2483);
    nor g2259(n2482 ,n2472 ,n2460);
    nor g2260(n2481 ,n2470 ,n2458);
    xnor g2261(n2480 ,n2446 ,n2283);
    xnor g2262(n2479 ,n2437 ,n2339);
    xnor g2263(n2478 ,n2431 ,n2327);
    xnor g2264(n2477 ,n2435 ,n2359);
    xnor g2265(n2476 ,n2439 ,n2343);
    nor g2266(n2483 ,n2441 ,n2465);
    not g2267(n2475 ,n2474);
    nor g2268(n2473 ,n2283 ,n2447);
    nor g2269(n2472 ,n2328 ,n2432);
    nor g2270(n2471 ,n2368 ,n2434);
    nor g2271(n2470 ,n2340 ,n2438);
    nor g2272(n2469 ,n2284 ,n2446);
    nor g2273(n2468 ,n2360 ,n2436);
    nor g2274(n2467 ,n2392 ,n2442);
    nor g2275(n2466 ,n2367 ,n2433);
    nor g2276(n2465 ,n2440 ,n2445);
    nor g2277(n2464 ,n2327 ,n2431);
    nor g2278(n2474 ,n2383 ,n2444);
    not g2279(n2462 ,n2461);
    not g2280(n2457 ,n2456);
    not g2281(n2455 ,n2454);
    not g2282(n2453 ,n2452);
    nor g2283(n2451 ,n2359 ,n2435);
    nor g2284(n2450 ,n2339 ,n2437);
    xnor g2285(n2449 ,n2415 ,n2357);
    xnor g2286(n2448 ,n2417 ,n2371);
    xnor g2287(n2463 ,n2414 ,n2350);
    xnor g2288(n2461 ,n2410 ,n2352);
    xnor g2289(n2460 ,n2407 ,n2379);
    xnor g2290(n2459 ,n2409 ,n2347);
    xnor g2291(n2458 ,n2408 ,n2351);
    xnor g2292(n2456 ,n2413 ,n2419);
    xnor g2293(n2454 ,n2412 ,n2393);
    xnor g2294(n2452 ,n2411 ,n2378);
    not g2295(n2447 ,n2446);
    nor g2296(n2445 ,n2358 ,n2415);
    nor g2297(n2444 ,n2399 ,n2420);
    nor g2298(n2443 ,n2371 ,n2418);
    nor g2299(n2442 ,n2372 ,n2417);
    nor g2300(n2441 ,n2357 ,n2416);
    nor g2301(n2446 ,n2396 ,n2427);
    not g2302(n2438 ,n2437);
    not g2303(n2436 ,n2435);
    not g2304(n2434 ,n2433);
    not g2305(n2432 ,n2431);
    xnor g2306(n2430 ,n2403 ,n2369);
    nor g2307(n2440 ,n2386 ,n2423);
    nor g2308(n2439 ,n2384 ,n2426);
    nor g2309(n2437 ,n2387 ,n2422);
    nor g2310(n2435 ,n2389 ,n2421);
    nor g2311(n2433 ,n2382 ,n2425);
    nor g2312(n2431 ,n2390 ,n2424);
    nor g2313(n2429 ,n2369 ,n2404);
    nor g2314(n2428 ,n2370 ,n2403);
    nor g2315(n2427 ,n2385 ,n2394);
    nor g2316(n2426 ,n2379 ,n2400);
    nor g2317(n2425 ,n2350 ,n2401);
    nor g2318(n2424 ,n2351 ,n2398);
    nor g2319(n2423 ,n2352 ,n2395);
    nor g2320(n2422 ,n2347 ,n2397);
    nor g2321(n2421 ,n2378 ,n2402);
    nor g2322(n3663 ,n2391 ,n2388);
    not g2323(n2420 ,n2419);
    not g2324(n2418 ,n2417);
    not g2325(n2416 ,n2415);
    xnor g2326(n2414 ,n2329 ,n2353);
    xnor g2327(n2413 ,n2335 ,n2361);
    xnor g2328(n2412 ,n2285 ,n2345);
    xnor g2329(n2411 ,n2365 ,n2333);
    xnor g2330(n2410 ,n2281 ,n2331);
    xnor g2331(n2409 ,n2337 ,n2375);
    xnor g2332(n2408 ,n2341 ,n2355);
    xnor g2333(n2407 ,n2373 ,n2363);
    xnor g2334(n2419 ,n2321 ,n2348);
    xnor g2335(n2417 ,n2323 ,n2377);
    xnor g2336(n2415 ,n2287 ,n2349);
    not g2337(n2406 ,n2405);
    not g2338(n2404 ,n2403);
    nor g2339(n2402 ,n2334 ,n2366);
    nor g2340(n2401 ,n2354 ,n2330);
    nor g2341(n2400 ,n2364 ,n2374);
    nor g2342(n2399 ,n2362 ,n2336);
    nor g2343(n2398 ,n2356 ,n2342);
    nor g2344(n2397 ,n2376 ,n2338);
    nor g2345(n2396 ,n2286 ,n2345);
    nor g2346(n2395 ,n2281 ,n2332);
    nor g2347(n2405 ,n2324 ,n2377);
    nor g2348(n2403 ,n2322 ,n2348);
    not g2349(n2394 ,n2393);
    not g2350(n2392 ,n2391);
    nor g2351(n2390 ,n2355 ,n2341);
    nor g2352(n2389 ,n2333 ,n2365);
    nor g2353(n2388 ,n2325 ,n2381);
    nor g2354(n2387 ,n2375 ,n2337);
    nor g2355(n2386 ,n2282 ,n2331);
    nor g2356(n2385 ,n2285 ,n2346);
    nor g2357(n2384 ,n2363 ,n2373);
    nor g2358(n2383 ,n2361 ,n2335);
    nor g2359(n2382 ,n2353 ,n2329);
    nor g2360(n2393 ,n2288 ,n2349);
    nor g2361(n2391 ,n2326 ,n2380);
    not g2362(n2381 ,n2380);
    not g2363(n2376 ,n2375);
    not g2364(n2374 ,n2373);
    not g2365(n2372 ,n2371);
    not g2366(n2370 ,n2369);
    not g2367(n2368 ,n2367);
    not g2368(n2366 ,n2365);
    not g2369(n2364 ,n2363);
    not g2370(n2362 ,n2361);
    not g2371(n2360 ,n2359);
    not g2372(n2358 ,n2357);
    not g2373(n2356 ,n2355);
    not g2374(n2354 ,n2353);
    nor g2375(n2380 ,n2250 ,n2299);
    nor g2376(n2379 ,n2257 ,n2316);
    nor g2377(n2378 ,n2270 ,n2318);
    nor g2378(n2377 ,n2266 ,n2311);
    nor g2379(n2375 ,n2245 ,n2294);
    nor g2380(n2373 ,n2276 ,n2306);
    nor g2381(n2371 ,n2251 ,n2290);
    nor g2382(n2369 ,n2279 ,n2292);
    nor g2383(n2367 ,n2260 ,n2314);
    nor g2384(n2365 ,n2275 ,n2302);
    nor g2385(n2363 ,n2249 ,n2289);
    nor g2386(n2361 ,n2268 ,n2315);
    nor g2387(n2359 ,n2252 ,n2300);
    nor g2388(n2357 ,n2269 ,n2301);
    nor g2389(n2355 ,n2254 ,n2313);
    nor g2390(n2353 ,n2267 ,n2298);
    not g2391(n2346 ,n2345);
    not g2392(n2344 ,n2343);
    not g2393(n2342 ,n2341);
    not g2394(n2340 ,n2339);
    not g2395(n2338 ,n2337);
    not g2396(n2336 ,n2335);
    not g2397(n2334 ,n2333);
    not g2398(n2332 ,n2331);
    not g2399(n2330 ,n2329);
    not g2400(n2328 ,n2327);
    nor g2401(n2352 ,n2278 ,n2312);
    nor g2402(n2351 ,n2246 ,n2296);
    nor g2403(n2350 ,n2256 ,n2307);
    nor g2404(n2349 ,n2280 ,n2305);
    nor g2405(n2348 ,n2248 ,n2317);
    nor g2406(n2347 ,n2277 ,n2310);
    nor g2407(n2345 ,n2258 ,n2319);
    nor g2408(n2343 ,n2247 ,n2320);
    nor g2409(n2341 ,n2272 ,n2303);
    nor g2410(n2339 ,n2273 ,n2295);
    nor g2411(n2337 ,n2265 ,n2293);
    nor g2412(n2335 ,n2255 ,n2308);
    nor g2413(n2333 ,n2274 ,n2304);
    nor g2414(n2331 ,n2259 ,n2291);
    nor g2415(n2329 ,n2253 ,n2309);
    nor g2416(n2327 ,n2271 ,n2297);
    not g2417(n2326 ,n2325);
    not g2418(n2324 ,n2323);
    not g2419(n2322 ,n2321);
    nor g2420(n2320 ,n2227 ,n2261);
    nor g2421(n2319 ,n2219 ,n2264);
    nor g2422(n2318 ,n2216 ,n2263);
    nor g2423(n2317 ,n2226 ,n2263);
    nor g2424(n2316 ,n2225 ,n2261);
    nor g2425(n2315 ,n2218 ,n2262);
    nor g2426(n2314 ,n2219 ,n2262);
    nor g2427(n2313 ,n2218 ,n2264);
    nor g2428(n2312 ,n2227 ,n2263);
    nor g2429(n2311 ,n2226 ,n2262);
    nor g2430(n2310 ,n2218 ,n2263);
    nor g2431(n2309 ,n2225 ,n2263);
    nor g2432(n2308 ,n2228 ,n2261);
    nor g2433(n2307 ,n2219 ,n2261);
    nor g2434(n2306 ,n2220 ,n2263);
    nor g2435(n2325 ,n2217 ,n2262);
    nor g2436(n2323 ,n2217 ,n2263);
    nor g2437(n2321 ,n2217 ,n2264);
    nor g2438(n2305 ,n2219 ,n2263);
    nor g2439(n2304 ,n2220 ,n2264);
    nor g2440(n2303 ,n2228 ,n2263);
    nor g2441(n2302 ,n2225 ,n2262);
    nor g2442(n2301 ,n2227 ,n2264);
    nor g2443(n2300 ,n2227 ,n2262);
    nor g2444(n3662 ,n2217 ,n2261);
    nor g2445(n2299 ,n2226 ,n2261);
    nor g2446(n2298 ,n2216 ,n2264);
    nor g2447(n2297 ,n2216 ,n2262);
    nor g2448(n2296 ,n2220 ,n2262);
    nor g2449(n2295 ,n2216 ,n2261);
    nor g2450(n2294 ,n2226 ,n2264);
    nor g2451(n2293 ,n2228 ,n2262);
    nor g2452(n2292 ,n2220 ,n2261);
    nor g2453(n2291 ,n2225 ,n2264);
    nor g2454(n2290 ,n2218 ,n2261);
    nor g2455(n2289 ,n2228 ,n2264);
    not g2456(n2288 ,n2287);
    not g2457(n2286 ,n2285);
    not g2458(n2284 ,n2283);
    not g2459(n2282 ,n2281);
    nor g2460(n2280 ,n2227 ,n2242);
    nor g2461(n2279 ,n2228 ,n2238);
    nor g2462(n2278 ,n2225 ,n2242);
    nor g2463(n2277 ,n2226 ,n2242);
    nor g2464(n2276 ,n2228 ,n2242);
    nor g2465(n2275 ,n2216 ,n2240);
    nor g2466(n2274 ,n2228 ,n2244);
    nor g2467(n2273 ,n2220 ,n2238);
    nor g2468(n2272 ,n2218 ,n2242);
    nor g2469(n2271 ,n2220 ,n2240);
    nor g2470(n2270 ,n2220 ,n2242);
    nor g2471(n2269 ,n2225 ,n2244);
    nor g2472(n2268 ,n2226 ,n2240);
    nor g2473(n2267 ,n2220 ,n2244);
    nor g2474(n2266 ,n2217 ,n2240);
    nor g2475(n2265 ,n2218 ,n2240);
    nor g2476(n2287 ,n2219 ,n2240);
    nor g2477(n2285 ,n2219 ,n2242);
    nor g2478(n2283 ,n2219 ,n2244);
    nor g2479(n2281 ,n2219 ,n2238);
    nor g2480(n2260 ,n2227 ,n2240);
    nor g2481(n2259 ,n2216 ,n2244);
    nor g2482(n2258 ,n2227 ,n2244);
    nor g2483(n2257 ,n2216 ,n2238);
    nor g2484(n2256 ,n2227 ,n2238);
    nor g2485(n2255 ,n2218 ,n2238);
    nor g2486(n2254 ,n2226 ,n2244);
    nor g2487(n2253 ,n2216 ,n2242);
    nor g2488(n2252 ,n2225 ,n2240);
    nor g2489(n2251 ,n2226 ,n2238);
    nor g2490(n2250 ,n2217 ,n2238);
    nor g2491(n2249 ,n2218 ,n2244);
    nor g2492(n2248 ,n2217 ,n2242);
    nor g2493(n2247 ,n2225 ,n2238);
    nor g2494(n2246 ,n2228 ,n2240);
    nor g2495(n2245 ,n2217 ,n2244);
    or g2496(n2264 ,n2243 ,n2233);
    or g2497(n2263 ,n2241 ,n2235);
    or g2498(n2262 ,n2239 ,n2236);
    or g2499(n2261 ,n2237 ,n2234);
    not g2500(n2244 ,n2243);
    nor g2501(n2243 ,n2230 ,n2221);
    not g2502(n2242 ,n2241);
    nor g2503(n2241 ,n2231 ,n2222);
    not g2504(n2240 ,n2239);
    nor g2505(n2239 ,n2232 ,n2224);
    not g2506(n2238 ,n2237);
    nor g2507(n2237 ,n2229 ,n2223);
    nor g2508(n2236 ,n28[1] ,n27[1]);
    nor g2509(n2235 ,n28[2] ,n27[2]);
    nor g2510(n2234 ,n28[0] ,n27[0]);
    nor g2511(n2233 ,n28[3] ,n27[3]);
    not g2512(n2232 ,n28[1]);
    not g2513(n2231 ,n28[2]);
    not g2514(n2230 ,n28[3]);
    not g2515(n2229 ,n28[0]);
    not g2516(n2228 ,n3679);
    not g2517(n2227 ,n3683);
    not g2518(n2226 ,n3677);
    not g2519(n2225 ,n3682);
    not g2520(n2224 ,n27[1]);
    not g2521(n2223 ,n27[0]);
    not g2522(n2222 ,n27[2]);
    not g2523(n2221 ,n27[3]);
    not g2524(n2220 ,n3680);
    not g2525(n2219 ,n3684);
    not g2526(n2218 ,n3678);
    not g2527(n2217 ,n3676);
    not g2528(n2216 ,n3681);
    or g2529(n30[11] ,n2766 ,n2851);
    xnor g2530(n30[10] ,n2774 ,n2850);
    nor g2531(n2851 ,n2769 ,n2850);
    nor g2532(n2850 ,n2793 ,n2849);
    xor g2533(n30[9] ,n2808 ,n2848);
    nor g2534(n2849 ,n2800 ,n2848);
    nor g2535(n2848 ,n2828 ,n2847);
    xnor g2536(n30[8] ,n2832 ,n2846);
    nor g2537(n2847 ,n2825 ,n2846);
    nor g2538(n2846 ,n2826 ,n2845);
    xnor g2539(n30[7] ,n2831 ,n2844);
    nor g2540(n2845 ,n2827 ,n2844);
    nor g2541(n2844 ,n2834 ,n2843);
    xor g2542(n30[6] ,n2839 ,n2842);
    nor g2543(n2843 ,n2837 ,n2842);
    nor g2544(n2842 ,n2833 ,n2841);
    xor g2545(n30[5] ,n2838 ,n2840);
    nor g2546(n2841 ,n2836 ,n2840);
    xnor g2547(n30[4] ,n2830 ,n2823);
    nor g2548(n2840 ,n2824 ,n2835);
    xnor g2549(n2839 ,n2819 ,n2821);
    xnor g2550(n2838 ,n2817 ,n2811);
    nor g2551(n2837 ,n2822 ,n2820);
    nor g2552(n2836 ,n2812 ,n2818);
    nor g2553(n2835 ,n2829 ,n2823);
    nor g2554(n2834 ,n2821 ,n2819);
    nor g2555(n2833 ,n2811 ,n2817);
    xnor g2556(n2832 ,n2795 ,n2814);
    xnor g2557(n2831 ,n2806 ,n2809);
    xnor g2558(n2830 ,n2803 ,n2786);
    xor g2559(n30[3] ,n2805 ,n2802);
    nor g2560(n2829 ,n2787 ,n2803);
    nor g2561(n2828 ,n2796 ,n2814);
    nor g2562(n2827 ,n2810 ,n2806);
    nor g2563(n2826 ,n2809 ,n2807);
    nor g2564(n2825 ,n2795 ,n2815);
    nor g2565(n2824 ,n2786 ,n2804);
    nor g2566(n2823 ,n2801 ,n2816);
    not g2567(n2822 ,n2821);
    nor g2568(n2821 ,n2799 ,n2813);
    not g2569(n2820 ,n2819);
    xnor g2570(n2819 ,n2789 ,n2779);
    not g2571(n2818 ,n2817);
    xnor g2572(n2817 ,n2790 ,n2775);
    nor g2573(n2816 ,n2802 ,n2797);
    not g2574(n2815 ,n2814);
    nor g2575(n2814 ,n2768 ,n2791);
    nor g2576(n2813 ,n2765 ,n2792);
    not g2577(n2812 ,n2811);
    nor g2578(n2811 ,n2751 ,n2794);
    not g2579(n2810 ,n2809);
    nor g2580(n2809 ,n2781 ,n2798);
    xnor g2581(n2808 ,n2784 ,n2736);
    not g2582(n2807 ,n2806);
    xnor g2583(n2806 ,n2773 ,n2788);
    xnor g2584(n2805 ,n2777 ,n2725);
    xor g2585(n30[2] ,n2772 ,n2729);
    not g2586(n2804 ,n2803);
    xnor g2587(n2803 ,n2758 ,n2780);
    nor g2588(n2801 ,n2726 ,n2778);
    nor g2589(n2800 ,n2737 ,n2785);
    nor g2590(n2799 ,n2741 ,n2776);
    nor g2591(n2798 ,n2783 ,n2779);
    nor g2592(n2797 ,n2725 ,n2777);
    nor g2593(n2802 ,n2771 ,n2782);
    not g2594(n2796 ,n2795);
    nor g2595(n2794 ,n2750 ,n2780);
    nor g2596(n2793 ,n2736 ,n2784);
    nor g2597(n2792 ,n2740 ,n2775);
    nor g2598(n2791 ,n2788 ,n2761);
    xor g2599(n2790 ,n2741 ,n2765);
    xnor g2600(n2789 ,n2763 ,n2685);
    xnor g2601(n2795 ,n2759 ,n2757);
    not g2602(n2787 ,n2786);
    not g2603(n2785 ,n2784);
    nor g2604(n2783 ,n2686 ,n2764);
    nor g2605(n2782 ,n2730 ,n2770);
    nor g2606(n2781 ,n2685 ,n2763);
    nor g2607(n2788 ,n2724 ,n2767);
    nor g2608(n2786 ,n2712 ,n2762);
    nor g2609(n2784 ,n2752 ,n2760);
    not g2610(n2778 ,n2777);
    not g2611(n2776 ,n2775);
    xnor g2612(n2774 ,n2755 ,n2581);
    xnor g2613(n2773 ,n2738 ,n2742);
    xnor g2614(n2772 ,n2734 ,n2705);
    xnor g2615(n2780 ,n2731 ,n2703);
    xnor g2616(n2779 ,n2732 ,n2746);
    xnor g2617(n2777 ,n2748 ,n2744);
    xnor g2618(n2775 ,n2733 ,n2674);
    nor g2619(n2771 ,n2705 ,n2735);
    nor g2620(n2770 ,n2706 ,n2734);
    nor g2621(n2769 ,n2581 ,n2756);
    nor g2622(n2768 ,n2739 ,n2742);
    nor g2623(n2767 ,n2714 ,n2747);
    nor g2624(n2766 ,n2582 ,n2755);
    not g2625(n2764 ,n2763);
    nor g2626(n2762 ,n2723 ,n2745);
    nor g2627(n2761 ,n2738 ,n2743);
    nor g2628(n2760 ,n2757 ,n2754);
    xnor g2629(n2759 ,n2719 ,n2701);
    xnor g2630(n2758 ,n2727 ,n2683);
    nor g2631(n2765 ,n2715 ,n2749);
    nor g2632(n2763 ,n2716 ,n2753);
    not g2633(n2756 ,n2755);
    nor g2634(n2754 ,n2702 ,n2719);
    nor g2635(n2753 ,n2675 ,n2721);
    nor g2636(n2752 ,n2701 ,n2720);
    nor g2637(n2751 ,n2683 ,n2728);
    nor g2638(n2750 ,n2684 ,n2727);
    nor g2639(n3639 ,n2729 ,n2717);
    nor g2640(n2749 ,n2691 ,n2722);
    xnor g2641(n2748 ,n2687 ,n2693);
    nor g2642(n2757 ,n2627 ,n2713);
    nor g2643(n2755 ,n2625 ,n2718);
    not g2644(n2747 ,n2746);
    not g2645(n2745 ,n2744);
    not g2646(n2743 ,n2742);
    not g2647(n2741 ,n2740);
    not g2648(n2739 ,n2738);
    not g2649(n2737 ,n2736);
    not g2650(n2735 ,n2734);
    xnor g2651(n2733 ,n2707 ,n2699);
    xnor g2652(n2732 ,n2583 ,n2695);
    xnor g2653(n2731 ,n2691 ,n2697);
    xnor g2654(n2746 ,n2682 ,n2597);
    xnor g2655(n2744 ,n2689 ,n2664);
    xnor g2656(n2742 ,n2654 ,n2692);
    xnor g2657(n2740 ,n2681 ,n2589);
    xnor g2658(n2738 ,n2680 ,n2591);
    xnor g2659(n2736 ,n2653 ,n2690);
    xnor g2660(n2734 ,n2709 ,n2676);
    not g2661(n2730 ,n2729);
    not g2662(n2728 ,n2727);
    not g2663(n2726 ,n2725);
    nor g2664(n2724 ,n2584 ,n2695);
    nor g2665(n2723 ,n2694 ,n2688);
    nor g2666(n2722 ,n2704 ,n2698);
    nor g2667(n2721 ,n2700 ,n2708);
    nor g2668(n2729 ,n2679 ,n2710);
    nor g2669(n2727 ,n2665 ,n2689);
    nor g2670(n2725 ,n2677 ,n2709);
    not g2671(n2720 ,n2719);
    nor g2672(n2718 ,n2620 ,n2690);
    nor g2673(n2717 ,n2678 ,n2711);
    nor g2674(n2716 ,n2699 ,n2707);
    nor g2675(n2715 ,n2703 ,n2697);
    nor g2676(n2714 ,n2583 ,n2696);
    nor g2677(n2713 ,n2618 ,n2692);
    nor g2678(n2712 ,n2693 ,n2687);
    xnor g2679(n2719 ,n2655 ,n2611);
    not g2680(n2711 ,n2710);
    not g2681(n2708 ,n2707);
    not g2682(n2706 ,n2705);
    not g2683(n2704 ,n2703);
    not g2684(n2702 ,n2701);
    not g2685(n2700 ,n2699);
    not g2686(n2698 ,n2697);
    not g2687(n2696 ,n2695);
    not g2688(n2694 ,n2693);
    nor g2689(n2710 ,n2641 ,n2661);
    nor g2690(n2709 ,n2643 ,n2670);
    nor g2691(n2707 ,n2639 ,n2669);
    nor g2692(n2705 ,n2634 ,n2668);
    nor g2693(n2703 ,n2644 ,n2666);
    nor g2694(n2701 ,n2617 ,n2663);
    nor g2695(n2699 ,n2642 ,n2673);
    nor g2696(n2697 ,n2637 ,n2667);
    nor g2697(n2695 ,n2640 ,n2671);
    nor g2698(n2693 ,n2633 ,n2660);
    not g2699(n2688 ,n2687);
    not g2700(n2686 ,n2685);
    not g2701(n2684 ,n2683);
    xnor g2702(n2682 ,n2651 ,n2587);
    xnor g2703(n2681 ,n2645 ,n2605);
    xnor g2704(n2680 ,n2649 ,n2607);
    nor g2705(n2692 ,n2622 ,n2658);
    xnor g2706(n2691 ,n2647 ,n2615);
    nor g2707(n2690 ,n2626 ,n2656);
    nor g2708(n2689 ,n2638 ,n2672);
    nor g2709(n2687 ,n2635 ,n2659);
    nor g2710(n2685 ,n2624 ,n2662);
    nor g2711(n2683 ,n2636 ,n2657);
    not g2712(n2679 ,n2678);
    not g2713(n2677 ,n2676);
    not g2714(n2675 ,n2674);
    nor g2715(n2673 ,n2573 ,n2630);
    nor g2716(n2672 ,n2574 ,n2629);
    nor g2717(n2671 ,n2574 ,n2630);
    nor g2718(n2670 ,n2566 ,n2631);
    nor g2719(n2669 ,n2574 ,n2632);
    nor g2720(n2668 ,n2573 ,n2629);
    nor g2721(n2667 ,n2574 ,n2631);
    nor g2722(n2666 ,n2573 ,n2632);
    nor g2723(n3638 ,n2565 ,n2629);
    nor g2724(n2678 ,n2565 ,n2631);
    nor g2725(n2676 ,n2565 ,n2632);
    nor g2726(n2674 ,n2616 ,n2648);
    not g2727(n2665 ,n2664);
    nor g2728(n2663 ,n2650 ,n2619);
    nor g2729(n2662 ,n2646 ,n2623);
    nor g2730(n2661 ,n2566 ,n2629);
    nor g2731(n2660 ,n2566 ,n2632);
    nor g2732(n2659 ,n2573 ,n2631);
    nor g2733(n2658 ,n2652 ,n2628);
    nor g2734(n2657 ,n2566 ,n2630);
    nor g2735(n2656 ,n2600 ,n2621);
    xnor g2736(n2655 ,n2609 ,n2599);
    xnor g2737(n2654 ,n2585 ,n2595);
    xnor g2738(n2653 ,n2613 ,n2593);
    nor g2739(n2664 ,n2565 ,n2630);
    not g2740(n2652 ,n2651);
    not g2741(n2650 ,n2649);
    not g2742(n2648 ,n2647);
    not g2743(n2646 ,n2645);
    nor g2744(n2644 ,n2566 ,n2604);
    nor g2745(n2643 ,n2565 ,n2602);
    nor g2746(n2642 ,n2566 ,n2601);
    nor g2747(n2641 ,n2565 ,n2603);
    nor g2748(n2640 ,n2573 ,n2601);
    nor g2749(n2639 ,n2573 ,n2604);
    nor g2750(n2638 ,n2573 ,n2603);
    nor g2751(n2637 ,n2573 ,n2602);
    nor g2752(n2636 ,n2565 ,n2601);
    nor g2753(n2635 ,n2566 ,n2602);
    nor g2754(n2634 ,n2566 ,n2603);
    nor g2755(n2633 ,n2565 ,n2604);
    nor g2756(n2651 ,n2574 ,n2604);
    nor g2757(n2649 ,n2574 ,n2601);
    nor g2758(n2647 ,n2574 ,n2603);
    nor g2759(n2645 ,n2574 ,n2602);
    nor g2760(n2628 ,n2587 ,n2597);
    nor g2761(n2627 ,n2596 ,n2586);
    nor g2762(n2626 ,n2612 ,n2610);
    nor g2763(n2625 ,n2594 ,n2614);
    nor g2764(n2624 ,n2606 ,n2590);
    nor g2765(n2623 ,n2605 ,n2589);
    nor g2766(n2622 ,n2588 ,n2598);
    nor g2767(n2621 ,n2611 ,n2609);
    nor g2768(n2620 ,n2593 ,n2613);
    nor g2769(n2619 ,n2607 ,n2591);
    nor g2770(n2618 ,n2595 ,n2585);
    nor g2771(n2617 ,n2608 ,n2592);
    xnor g2772(n2632 ,n3647 ,n4[2]);
    xnor g2773(n2631 ,n3646 ,n4[1]);
    xnor g2774(n2630 ,n3648 ,n4[3]);
    xnor g2775(n2629 ,n3645 ,n4[0]);
    not g2776(n2616 ,n2615);
    not g2777(n2614 ,n2613);
    not g2778(n2612 ,n2611);
    not g2779(n2610 ,n2609);
    not g2780(n2608 ,n2607);
    not g2781(n2606 ,n2605);
    nor g2782(n2615 ,n2565 ,n2575);
    nor g2783(n2613 ,n2574 ,n2567);
    nor g2784(n2611 ,n2573 ,n2567);
    nor g2785(n2609 ,n2574 ,n2569);
    nor g2786(n2607 ,n2565 ,n2568);
    nor g2787(n2605 ,n2565 ,n2569);
    or g2788(n2604 ,n2571 ,n2580);
    or g2789(n2603 ,n2579 ,n2578);
    or g2790(n2602 ,n2570 ,n2576);
    or g2791(n2601 ,n2577 ,n2572);
    not g2792(n2600 ,n2599);
    not g2793(n2598 ,n2597);
    not g2794(n2596 ,n2595);
    not g2795(n2594 ,n2593);
    not g2796(n2592 ,n2591);
    not g2797(n2590 ,n2589);
    not g2798(n2588 ,n2587);
    not g2799(n2586 ,n2585);
    not g2800(n2584 ,n2583);
    not g2801(n2582 ,n2581);
    nor g2802(n2599 ,n2566 ,n2568);
    nor g2803(n2597 ,n2573 ,n2575);
    nor g2804(n2595 ,n2566 ,n2567);
    nor g2805(n2593 ,n2573 ,n2568);
    nor g2806(n2591 ,n2574 ,n2575);
    nor g2807(n2589 ,n2566 ,n2575);
    nor g2808(n2587 ,n2565 ,n2567);
    nor g2809(n2585 ,n2573 ,n2569);
    nor g2810(n2583 ,n2566 ,n2569);
    nor g2811(n2581 ,n2574 ,n2568);
    not g2812(n2580 ,n4[2]);
    not g2813(n2579 ,n3645);
    not g2814(n2578 ,n4[0]);
    not g2815(n2577 ,n3648);
    not g2816(n2576 ,n4[1]);
    not g2817(n2575 ,n4[4]);
    not g2818(n2574 ,n5[3]);
    not g2819(n2573 ,n5[2]);
    not g2820(n2572 ,n4[3]);
    not g2821(n2571 ,n3647);
    not g2822(n2570 ,n3646);
    not g2823(n2569 ,n4[5]);
    not g2824(n2568 ,n4[7]);
    not g2825(n2567 ,n4[6]);
    not g2826(n2566 ,n5[1]);
    not g2827(n2565 ,n5[0]);
    or g2828(n3661 ,n3300 ,n3368);
    xor g2829(n3660 ,n3308 ,n3367);
    nor g2830(n3368 ,n3301 ,n3367);
    nor g2831(n3367 ,n3332 ,n3366);
    xnor g2832(n3659 ,n3342 ,n3365);
    nor g2833(n3366 ,n3333 ,n3365);
    nor g2834(n3365 ,n3345 ,n3364);
    xor g2835(n3658 ,n3349 ,n3363);
    nor g2836(n3364 ,n3346 ,n3363);
    nor g2837(n3363 ,n3350 ,n3362);
    xor g2838(n3657 ,n3356 ,n3361);
    nor g2839(n3362 ,n3354 ,n3361);
    nor g2840(n3361 ,n3352 ,n3360);
    xor g2841(n3656 ,n3355 ,n3359);
    nor g2842(n3360 ,n3353 ,n3359);
    nor g2843(n3359 ,n3344 ,n3358);
    xor g2844(n3655 ,n3348 ,n3357);
    nor g2845(n3358 ,n3347 ,n3357);
    nor g2846(n3357 ,n3334 ,n3351);
    xnor g2847(n3356 ,n3339 ,n3329);
    xnor g2848(n3355 ,n3337 ,n3335);
    xnor g2849(n3654 ,n3341 ,n3343);
    nor g2850(n3354 ,n3330 ,n3340);
    nor g2851(n3353 ,n3336 ,n3338);
    nor g2852(n3352 ,n3335 ,n3337);
    nor g2853(n3351 ,n3331 ,n3343);
    nor g2854(n3350 ,n3329 ,n3339);
    xnor g2855(n3349 ,n3310 ,n3327);
    xnor g2856(n3348 ,n3325 ,n3321);
    xnor g2857(n3653 ,n3323 ,n3314);
    nor g2858(n3347 ,n3322 ,n3326);
    nor g2859(n3346 ,n3328 ,n3311);
    nor g2860(n3345 ,n3327 ,n3310);
    nor g2861(n3344 ,n3321 ,n3325);
    nor g2862(n3343 ,n3317 ,n3324);
    xnor g2863(n3342 ,n3276 ,n3319);
    xnor g2864(n3341 ,n3312 ,n3294);
    not g2865(n3340 ,n3339);
    xnor g2866(n3339 ,n3307 ,n3287);
    not g2867(n3338 ,n3337);
    xnor g2868(n3337 ,n3306 ,n3268);
    not g2869(n3336 ,n3335);
    nor g2870(n3334 ,n3294 ,n3313);
    nor g2871(n3333 ,n3276 ,n3320);
    nor g2872(n3332 ,n3277 ,n3319);
    nor g2873(n3331 ,n3295 ,n3312);
    nor g2874(n3335 ,n3299 ,n3316);
    not g2875(n3330 ,n3329);
    not g2876(n3328 ,n3327);
    not g2877(n3326 ,n3325);
    nor g2878(n3324 ,n3314 ,n3318);
    xnor g2879(n3652 ,n3289 ,n3288);
    xnor g2880(n3323 ,n3296 ,n3266);
    nor g2881(n3329 ,n3293 ,n3309);
    nor g2882(n3327 ,n3303 ,n3315);
    xnor g2883(n3325 ,n3290 ,n3274);
    not g2884(n3322 ,n3321);
    not g2885(n3320 ,n3319);
    nor g2886(n3318 ,n3267 ,n3296);
    nor g2887(n3317 ,n3266 ,n3297);
    nor g2888(n3316 ,n3237 ,n3302);
    nor g2889(n3315 ,n3287 ,n3291);
    nor g2890(n3321 ,n3282 ,n3298);
    nor g2891(n3319 ,n3260 ,n3292);
    not g2892(n3313 ,n3312);
    not g2893(n3311 ,n3310);
    nor g2894(n3309 ,n3268 ,n3304);
    xnor g2895(n3308 ,n3285 ,n3094);
    xnor g2896(n3307 ,n3232 ,n3278);
    xnor g2897(n3306 ,n3253 ,n3272);
    nor g2898(n3314 ,n3284 ,n3305);
    xnor g2899(n3312 ,n3270 ,n3255);
    xnor g2900(n3310 ,n3269 ,n3280);
    nor g2901(n3305 ,n3288 ,n3281);
    nor g2902(n3304 ,n3254 ,n3273);
    nor g2903(n3303 ,n3233 ,n3279);
    nor g2904(n3302 ,n3252 ,n3275);
    nor g2905(n3301 ,n3095 ,n3286);
    nor g2906(n3300 ,n3094 ,n3285);
    nor g2907(n3299 ,n3251 ,n3274);
    nor g2908(n3298 ,n3238 ,n3283);
    not g2909(n3297 ,n3296);
    not g2910(n3295 ,n3294);
    nor g2911(n3293 ,n3253 ,n3272);
    nor g2912(n3292 ,n3280 ,n3261);
    nor g2913(n3291 ,n3232 ,n3278);
    xor g2914(n3651 ,n3249 ,n3225);
    xnor g2915(n3290 ,n3251 ,n3237);
    xnor g2916(n3289 ,n3257 ,n3173);
    xnor g2917(n3296 ,n3250 ,n3259);
    nor g2918(n3294 ,n3240 ,n3271);
    not g2919(n3286 ,n3285);
    nor g2920(n3284 ,n3173 ,n3258);
    nor g2921(n3283 ,n3230 ,n3256);
    nor g2922(n3282 ,n3231 ,n3255);
    nor g2923(n3281 ,n3174 ,n3257);
    nor g2924(n3288 ,n3239 ,n3263);
    nor g2925(n3287 ,n3218 ,n3264);
    nor g2926(n3285 ,n3192 ,n3265);
    not g2927(n3279 ,n3278);
    not g2928(n3277 ,n3276);
    not g2929(n3275 ,n3274);
    not g2930(n3273 ,n3272);
    nor g2931(n3271 ,n3243 ,n3259);
    xnor g2932(n3270 ,n3230 ,n3238);
    xnor g2933(n3269 ,n3234 ,n3245);
    nor g2934(n3280 ,n3223 ,n3262);
    xnor g2935(n3278 ,n3228 ,n3247);
    xnor g2936(n3276 ,n3203 ,n3248);
    xnor g2937(n3274 ,n3227 ,n3226);
    xnor g2938(n3272 ,n3229 ,n3236);
    not g2939(n3267 ,n3266);
    nor g2940(n3265 ,n3190 ,n3248);
    nor g2941(n3264 ,n3224 ,n3236);
    nor g2942(n3263 ,n3225 ,n3244);
    nor g2943(n3262 ,n3222 ,n3247);
    nor g2944(n3261 ,n3246 ,n3235);
    nor g2945(n3260 ,n3245 ,n3234);
    nor g2946(n3268 ,n3221 ,n3241);
    nor g2947(n3266 ,n3194 ,n3242);
    not g2948(n3258 ,n3257);
    not g2949(n3256 ,n3255);
    not g2950(n3254 ,n3253);
    not g2951(n3252 ,n3251);
    xnor g2952(n3650 ,n3038 ,n3202);
    xnor g2953(n3250 ,n3211 ,n3179);
    xnor g2954(n3249 ,n3154 ,n3209);
    xnor g2955(n3259 ,n3205 ,n3142);
    xnor g2956(n3257 ,n3206 ,n3213);
    xnor g2957(n3255 ,n3200 ,n3185);
    xnor g2958(n3253 ,n3204 ,n3160);
    xnor g2959(n3251 ,n3201 ,n3134);
    not g2960(n3246 ,n3245);
    nor g2961(n3244 ,n3154 ,n3209);
    nor g2962(n3243 ,n3180 ,n3211);
    nor g2963(n3242 ,n3169 ,n3214);
    nor g2964(n3241 ,n3220 ,n3226);
    nor g2965(n3240 ,n3179 ,n3212);
    nor g2966(n3239 ,n3155 ,n3210);
    nor g2967(n3248 ,n3187 ,n3215);
    nor g2968(n3247 ,n3198 ,n3217);
    nor g2969(n3245 ,n3189 ,n3207);
    not g2970(n3235 ,n3234);
    not g2971(n3233 ,n3232);
    not g2972(n3231 ,n3230);
    xnor g2973(n3229 ,n3177 ,n3175);
    xnor g2974(n3228 ,n3124 ,n3181);
    xnor g2975(n3227 ,n3183 ,n3096);
    nor g2976(n3238 ,n3196 ,n3216);
    nor g2977(n3237 ,n3197 ,n3219);
    nor g2978(n3236 ,n3195 ,n3208);
    xnor g2979(n3234 ,n3166 ,n3140);
    xnor g2980(n3232 ,n3168 ,n3132);
    xnor g2981(n3230 ,n3167 ,n3162);
    nor g2982(n3224 ,n3176 ,n3178);
    nor g2983(n3223 ,n3181 ,n3125);
    nor g2984(n3222 ,n3182 ,n3124);
    nor g2985(n3221 ,n3096 ,n3183);
    nor g2986(n3220 ,n3097 ,n3184);
    nor g2987(n3219 ,n3185 ,n3170);
    nor g2988(n3218 ,n3175 ,n3177);
    nor g2989(n3217 ,n3119 ,n3199);
    nor g2990(n3216 ,n3106 ,n3171);
    nor g2991(n3215 ,n3102 ,n3186);
    nor g2992(n3226 ,n3153 ,n3191);
    nor g2993(n3225 ,n3073 ,n3193);
    not g2994(n3214 ,n3213);
    not g2995(n3212 ,n3211);
    not g2996(n3210 ,n3209);
    nor g2997(n3208 ,n3101 ,n3172);
    nor g2998(n3207 ,n3103 ,n3188);
    xnor g2999(n3206 ,n3130 ,n3128);
    xnor g3000(n3205 ,n3138 ,n3106);
    xnor g3001(n3204 ,n3156 ,n3119);
    xnor g3002(n3203 ,n3144 ,n3158);
    xnor g3003(n3202 ,n3164 ,n2882);
    xnor g3004(n3201 ,n3136 ,n3101);
    xnor g3005(n3200 ,n3122 ,n3126);
    xnor g3006(n3213 ,n3120 ,n3100);
    xnor g3007(n3211 ,n3121 ,n3105);
    xnor g3008(n3209 ,n3146 ,n3118);
    nor g3009(n3199 ,n3156 ,n3160);
    nor g3010(n3198 ,n3157 ,n3161);
    nor g3011(n3197 ,n3123 ,n3127);
    nor g3012(n3196 ,n3143 ,n3139);
    nor g3013(n3195 ,n3137 ,n3135);
    nor g3014(n3194 ,n3131 ,n3129);
    nor g3015(n3193 ,n3074 ,n3165);
    nor g3016(n3192 ,n3158 ,n3145);
    nor g3017(n3191 ,n3163 ,n3147);
    nor g3018(n3190 ,n3159 ,n3144);
    nor g3019(n3189 ,n3098 ,n3133);
    nor g3020(n3188 ,n3099 ,n3132);
    nor g3021(n3187 ,n3092 ,n3140);
    nor g3022(n3186 ,n3093 ,n3141);
    not g3023(n3184 ,n3183);
    not g3024(n3182 ,n3181);
    not g3025(n3180 ,n3179);
    not g3026(n3178 ,n3177);
    not g3027(n3176 ,n3175);
    not g3028(n3174 ,n3173);
    nor g3029(n3172 ,n3136 ,n3134);
    nor g3030(n3171 ,n3142 ,n3138);
    nor g3031(n3170 ,n3122 ,n3126);
    nor g3032(n3169 ,n3130 ,n3128);
    xnor g3033(n3168 ,n3103 ,n3098);
    xnor g3034(n3167 ,n3115 ,n3113);
    xnor g3035(n3166 ,n3102 ,n3092);
    nor g3036(n3185 ,n3111 ,n3152);
    xnor g3037(n3183 ,n3059 ,n3104);
    nor g3038(n3181 ,n3030 ,n3151);
    nor g3039(n3179 ,n3108 ,n3148);
    xnor g3040(n3177 ,n3053 ,n3117);
    nor g3041(n3175 ,n3023 ,n3150);
    nor g3042(n3173 ,n3112 ,n3149);
    not g3043(n3165 ,n3164);
    not g3044(n3163 ,n3162);
    not g3045(n3161 ,n3160);
    not g3046(n3159 ,n3158);
    not g3047(n3157 ,n3156);
    not g3048(n3155 ,n3154);
    nor g3049(n3153 ,n3113 ,n3115);
    nor g3050(n3152 ,n3105 ,n3110);
    nor g3051(n3151 ,n3013 ,n3117);
    nor g3052(n3150 ,n2999 ,n3104);
    nor g3053(n3149 ,n3118 ,n3109);
    nor g3054(n3148 ,n3100 ,n3107);
    nor g3055(n3147 ,n3114 ,n3116);
    xnor g3056(n3146 ,n3068 ,n2884);
    xnor g3057(n3164 ,n3061 ,n2902);
    xnor g3058(n3162 ,n3060 ,n2930);
    xnor g3059(n3160 ,n3063 ,n2888);
    nor g3060(n3158 ,n3026 ,n3091);
    xnor g3061(n3156 ,n3048 ,n2993);
    xnor g3062(n3154 ,n3071 ,n2948);
    not g3063(n3145 ,n3144);
    not g3064(n3143 ,n3142);
    not g3065(n3141 ,n3140);
    not g3066(n3139 ,n3138);
    not g3067(n3137 ,n3136);
    not g3068(n3135 ,n3134);
    not g3069(n3133 ,n3132);
    not g3070(n3131 ,n3130);
    not g3071(n3129 ,n3128);
    not g3072(n3127 ,n3126);
    not g3073(n3125 ,n3124);
    not g3074(n3123 ,n3122);
    xnor g3075(n3121 ,n3064 ,n3041);
    xnor g3076(n3120 ,n3066 ,n3039);
    xnor g3077(n3144 ,n3049 ,n3045);
    xnor g3078(n3142 ,n3055 ,n2921);
    xnor g3079(n3140 ,n3050 ,n3070);
    xnor g3080(n3138 ,n3054 ,n2944);
    xnor g3081(n3136 ,n3052 ,n2981);
    xnor g3082(n3134 ,n3062 ,n2900);
    xnor g3083(n3132 ,n3072 ,n2983);
    xnor g3084(n3130 ,n3047 ,n2978);
    xnor g3085(n3128 ,n3058 ,n2964);
    xnor g3086(n3126 ,n3056 ,n3043);
    xnor g3087(n3124 ,n3057 ,n2991);
    xnor g3088(n3122 ,n3051 ,n2958);
    not g3089(n3116 ,n3115);
    not g3090(n3114 ,n3113);
    nor g3091(n3112 ,n2885 ,n3068);
    nor g3092(n3111 ,n3042 ,n3064);
    nor g3093(n3110 ,n3041 ,n3065);
    nor g3094(n3109 ,n2884 ,n3069);
    nor g3095(n3108 ,n3040 ,n3066);
    nor g3096(n3107 ,n3039 ,n3067);
    nor g3097(n3119 ,n3024 ,n3086);
    nor g3098(n3118 ,n3018 ,n3075);
    nor g3099(n3117 ,n3032 ,n3079);
    nor g3100(n3115 ,n3034 ,n3088);
    nor g3101(n3113 ,n3035 ,n3080);
    not g3102(n3099 ,n3098);
    not g3103(n3097 ,n3096);
    not g3104(n3095 ,n3094);
    not g3105(n3093 ,n3092);
    nor g3106(n3091 ,n3006 ,n3070);
    nor g3107(n3106 ,n3021 ,n3077);
    nor g3108(n3105 ,n3036 ,n3082);
    nor g3109(n3104 ,n3020 ,n3078);
    nor g3110(n3103 ,n3008 ,n3089);
    nor g3111(n3102 ,n3025 ,n3087);
    nor g3112(n3101 ,n3027 ,n3085);
    nor g3113(n3100 ,n3022 ,n3076);
    nor g3114(n3098 ,n3029 ,n3083);
    nor g3115(n3096 ,n3033 ,n3081);
    nor g3116(n3094 ,n3031 ,n3084);
    nor g3117(n3092 ,n3028 ,n3090);
    nor g3118(n3090 ,n2984 ,n3005);
    nor g3119(n3089 ,n2918 ,n3011);
    nor g3120(n3088 ,n2922 ,n3002);
    nor g3121(n3087 ,n2992 ,n3014);
    nor g3122(n3086 ,n2997 ,n3010);
    nor g3123(n3085 ,n2980 ,n3012);
    nor g3124(n3084 ,n3004 ,n3046);
    nor g3125(n3083 ,n2994 ,n3003);
    nor g3126(n3082 ,n2979 ,n3007);
    nor g3127(n3081 ,n3009 ,n3044);
    nor g3128(n3080 ,n2927 ,n3001);
    nor g3129(n3079 ,n2982 ,n3016);
    nor g3130(n3078 ,n2931 ,n3019);
    nor g3131(n3077 ,n2985 ,n3000);
    nor g3132(n3076 ,n2924 ,n3017);
    nor g3133(n3075 ,n2990 ,n2998);
    nor g3134(n3074 ,n2882 ,n3038);
    nor g3135(n3649 ,n3015 ,n3038);
    nor g3136(n3073 ,n2883 ,n3037);
    xnor g3137(n3072 ,n2976 ,n2908);
    xnor g3138(n3071 ,n2923 ,n2890);
    not g3139(n3069 ,n3068);
    not g3140(n3067 ,n3066);
    not g3141(n3065 ,n3064);
    xor g3142(n3063 ,n2918 ,n2972);
    xor g3143(n3062 ,n2997 ,n2966);
    xor g3144(n3061 ,n2990 ,n2912);
    xnor g3145(n3060 ,n2876 ,n2896);
    xnor g3146(n3059 ,n2914 ,n2946);
    xor g3147(n3058 ,n2985 ,n2894);
    xnor g3148(n3057 ,n2878 ,n2942);
    xnor g3149(n3056 ,n2910 ,n2962);
    xnor g3150(n3055 ,n2906 ,n2886);
    xor g3151(n3054 ,n2927 ,n2954);
    xnor g3152(n3053 ,n2898 ,n2960);
    xnor g3153(n3052 ,n2880 ,n2970);
    xor g3154(n3051 ,n2980 ,n2904);
    xnor g3155(n3050 ,n2940 ,n2892);
    xnor g3156(n3049 ,n2968 ,n2938);
    xnor g3157(n3048 ,n2974 ,n2950);
    xnor g3158(n3047 ,n2952 ,n2956);
    xnor g3159(n3070 ,n2925 ,n2932);
    xnor g3160(n3068 ,n2995 ,n2916);
    xnor g3161(n3066 ,n2988 ,n2928);
    xnor g3162(n3064 ,n2986 ,n2919);
    not g3163(n3046 ,n3045);
    not g3164(n3044 ,n3043);
    not g3165(n3042 ,n3041);
    not g3166(n3040 ,n3039);
    not g3167(n3037 ,n3038);
    nor g3168(n3036 ,n2957 ,n2953);
    nor g3169(n3035 ,n2955 ,n2945);
    nor g3170(n3034 ,n2887 ,n2907);
    nor g3171(n3033 ,n2963 ,n2911);
    nor g3172(n3032 ,n2971 ,n2881);
    nor g3173(n3031 ,n2939 ,n2969);
    nor g3174(n3030 ,n2961 ,n2899);
    nor g3175(n3029 ,n2951 ,n2975);
    nor g3176(n3028 ,n2909 ,n2977);
    nor g3177(n3027 ,n2959 ,n2905);
    nor g3178(n3026 ,n2893 ,n2941);
    nor g3179(n3025 ,n2943 ,n2879);
    nor g3180(n3024 ,n2901 ,n2967);
    nor g3181(n3023 ,n2947 ,n2915);
    nor g3182(n3022 ,n2891 ,n2949);
    nor g3183(n3021 ,n2895 ,n2965);
    nor g3184(n3020 ,n2897 ,n2877);
    nor g3185(n3045 ,n2933 ,n2926);
    nor g3186(n3043 ,n2920 ,n2987);
    nor g3187(n3041 ,n2929 ,n2989);
    nor g3188(n3039 ,n2917 ,n2996);
    nor g3189(n3038 ,n2937 ,n2935);
    nor g3190(n3019 ,n2896 ,n2876);
    nor g3191(n3018 ,n2913 ,n2903);
    nor g3192(n3017 ,n2890 ,n2948);
    nor g3193(n3016 ,n2970 ,n2880);
    nor g3194(n3015 ,n2936 ,n2934);
    nor g3195(n3014 ,n2942 ,n2878);
    nor g3196(n3013 ,n2960 ,n2898);
    nor g3197(n3012 ,n2958 ,n2904);
    nor g3198(n3011 ,n2888 ,n2972);
    nor g3199(n3010 ,n2900 ,n2966);
    nor g3200(n3009 ,n2962 ,n2910);
    nor g3201(n3008 ,n2889 ,n2973);
    nor g3202(n3007 ,n2956 ,n2952);
    nor g3203(n3006 ,n2892 ,n2940);
    nor g3204(n3005 ,n2908 ,n2976);
    nor g3205(n3004 ,n2938 ,n2968);
    nor g3206(n3003 ,n2950 ,n2974);
    nor g3207(n3002 ,n2886 ,n2906);
    nor g3208(n3001 ,n2954 ,n2944);
    nor g3209(n3000 ,n2894 ,n2964);
    nor g3210(n2999 ,n2946 ,n2914);
    nor g3211(n2998 ,n2912 ,n2902);
    not g3212(n2996 ,n2995);
    not g3213(n2994 ,n2993);
    not g3214(n2992 ,n2991);
    not g3215(n2989 ,n2988);
    not g3216(n2987 ,n2986);
    not g3217(n2984 ,n2983);
    not g3218(n2982 ,n2981);
    not g3219(n2979 ,n2978);
    not g3220(n2977 ,n2976);
    not g3221(n2975 ,n2974);
    not g3222(n2973 ,n2972);
    not g3223(n2971 ,n2970);
    not g3224(n2969 ,n2968);
    not g3225(n2967 ,n2966);
    not g3226(n2965 ,n2964);
    not g3227(n2963 ,n2962);
    not g3228(n2961 ,n2960);
    not g3229(n2959 ,n2958);
    not g3230(n2957 ,n2956);
    not g3231(n2955 ,n2954);
    not g3232(n2953 ,n2952);
    not g3233(n2951 ,n2950);
    not g3234(n2949 ,n2948);
    not g3235(n2947 ,n2946);
    not g3236(n2945 ,n2944);
    not g3237(n2943 ,n2942);
    not g3238(n2941 ,n2940);
    not g3239(n2939 ,n2938);
    or g3240(n2997 ,n2852 ,n2868);
    nor g3241(n2995 ,n2856 ,n2857);
    nor g3242(n2993 ,n2854 ,n2859);
    nor g3243(n2991 ,n2852 ,n2863);
    or g3244(n2990 ,n2865 ,n2874);
    nor g3245(n2988 ,n2856 ,n2860);
    nor g3246(n2986 ,n2856 ,n2870);
    or g3247(n2985 ,n2852 ,n2874);
    nor g3248(n2983 ,n2865 ,n2861);
    nor g3249(n2981 ,n2854 ,n2870);
    or g3250(n2980 ,n2852 ,n2875);
    nor g3251(n2978 ,n2866 ,n2869);
    nor g3252(n2976 ,n2853 ,n2862);
    nor g3253(n2974 ,n2856 ,n2862);
    nor g3254(n2972 ,n2855 ,n2861);
    nor g3255(n2970 ,n2864 ,n2862);
    nor g3256(n2968 ,n2852 ,n2861);
    nor g3257(n2966 ,n2855 ,n2873);
    nor g3258(n2964 ,n2855 ,n2868);
    nor g3259(n2962 ,n2865 ,n2858);
    nor g3260(n2960 ,n2865 ,n2873);
    nor g3261(n2958 ,n2853 ,n2870);
    nor g3262(n2956 ,n2853 ,n2857);
    nor g3263(n2954 ,n2854 ,n2857);
    nor g3264(n2952 ,n2865 ,n2875);
    nor g3265(n2950 ,n2864 ,n2872);
    nor g3266(n2948 ,n2865 ,n2869);
    nor g3267(n2946 ,n2865 ,n2863);
    nor g3268(n2944 ,n2855 ,n2858);
    nor g3269(n2942 ,n2854 ,n2867);
    nor g3270(n2940 ,n2852 ,n2873);
    nor g3271(n2938 ,n2854 ,n2872);
    not g3272(n2937 ,n2936);
    not g3273(n2935 ,n2934);
    not g3274(n2933 ,n2932);
    not g3275(n2931 ,n2930);
    not g3276(n2929 ,n2928);
    not g3277(n2926 ,n2925);
    not g3278(n2924 ,n2923);
    not g3279(n2922 ,n2921);
    not g3280(n2920 ,n2919);
    not g3281(n2917 ,n2916);
    not g3282(n2915 ,n2914);
    not g3283(n2913 ,n2912);
    not g3284(n2911 ,n2910);
    not g3285(n2909 ,n2908);
    not g3286(n2907 ,n2906);
    not g3287(n2905 ,n2904);
    not g3288(n2903 ,n2902);
    not g3289(n2901 ,n2900);
    not g3290(n2899 ,n2898);
    not g3291(n2897 ,n2896);
    not g3292(n2895 ,n2894);
    not g3293(n2893 ,n2892);
    not g3294(n2891 ,n2890);
    not g3295(n2889 ,n2888);
    not g3296(n2887 ,n2886);
    not g3297(n2885 ,n2884);
    not g3298(n2883 ,n2882);
    not g3299(n2881 ,n2880);
    not g3300(n2879 ,n2878);
    not g3301(n2877 ,n2876);
    nor g3302(n2936 ,n2864 ,n2871);
    nor g3303(n2934 ,n2855 ,n2874);
    nor g3304(n2932 ,n2853 ,n2872);
    nor g3305(n2930 ,n2854 ,n2860);
    nor g3306(n2928 ,n2864 ,n2870);
    or g3307(n2927 ,n2852 ,n2869);
    nor g3308(n2925 ,n2854 ,n2862);
    nor g3309(n2923 ,n2866 ,n2874);
    nor g3310(n2921 ,n2866 ,n2875);
    nor g3311(n2919 ,n2864 ,n2859);
    or g3312(n2918 ,n2852 ,n2858);
    nor g3313(n2916 ,n2864 ,n2860);
    nor g3314(n2914 ,n2866 ,n2858);
    nor g3315(n2912 ,n2864 ,n2857);
    nor g3316(n2910 ,n2866 ,n2868);
    nor g3317(n2908 ,n2856 ,n2872);
    nor g3318(n2906 ,n2865 ,n2868);
    nor g3319(n2904 ,n2855 ,n2863);
    nor g3320(n2902 ,n2855 ,n2869);
    nor g3321(n2900 ,n2853 ,n2859);
    nor g3322(n2898 ,n2866 ,n2863);
    nor g3323(n2896 ,n2864 ,n2867);
    nor g3324(n2894 ,n2854 ,n2871);
    nor g3325(n2892 ,n2866 ,n2861);
    nor g3326(n2890 ,n2855 ,n2875);
    nor g3327(n2888 ,n2853 ,n2867);
    nor g3328(n2886 ,n2853 ,n2860);
    nor g3329(n2884 ,n2853 ,n2871);
    nor g3330(n2882 ,n2856 ,n2871);
    nor g3331(n2880 ,n2856 ,n2867);
    nor g3332(n2878 ,n2866 ,n2873);
    nor g3333(n2876 ,n2856 ,n2859);
    not g3334(n2875 ,n4[2]);
    not g3335(n2874 ,n4[0]);
    not g3336(n2873 ,n4[6]);
    not g3337(n2872 ,n26[7]);
    not g3338(n2871 ,n26[0]);
    not g3339(n2870 ,n26[3]);
    not g3340(n2869 ,n4[1]);
    not g3341(n2868 ,n4[3]);
    not g3342(n2867 ,n26[5]);
    not g3343(n2866 ,n27[2]);
    not g3344(n2865 ,n27[1]);
    not g3345(n2864 ,n28[0]);
    not g3346(n2863 ,n4[5]);
    not g3347(n2862 ,n26[6]);
    not g3348(n2861 ,n4[7]);
    not g3349(n2860 ,n26[2]);
    not g3350(n2859 ,n26[4]);
    not g3351(n2858 ,n4[4]);
    not g3352(n2857 ,n26[1]);
    not g3353(n2856 ,n28[1]);
    not g3354(n2855 ,n27[0]);
    not g3355(n2854 ,n28[3]);
    not g3356(n2853 ,n28[2]);
    not g3357(n2852 ,n27[3]);
    nor g3358(n3684 ,n3380 ,n3409);
    xnor g3359(n3683 ,n3388 ,n3408);
    nor g3360(n3409 ,n3388 ,n3408);
    nor g3361(n3408 ,n3381 ,n3407);
    xor g3362(n3682 ,n3389 ,n3405);
    nor g3363(n3407 ,n3389 ,n3406);
    not g3364(n3406 ,n3405);
    nor g3365(n3405 ,n3387 ,n3404);
    xor g3366(n3681 ,n3392 ,n3403);
    nor g3367(n3404 ,n3392 ,n3403);
    nor g3368(n3403 ,n3385 ,n3402);
    xor g3369(n3680 ,n3391 ,n3401);
    nor g3370(n3402 ,n3391 ,n3401);
    nor g3371(n3401 ,n3383 ,n3400);
    xor g3372(n3679 ,n3394 ,n3399);
    nor g3373(n3400 ,n3394 ,n3399);
    nor g3374(n3399 ,n3386 ,n3398);
    xnor g3375(n3678 ,n3393 ,n3396);
    nor g3376(n3398 ,n3393 ,n3397);
    not g3377(n3397 ,n3396);
    nor g3378(n3396 ,n3379 ,n3395);
    xnor g3379(n3677 ,n3390 ,n3384);
    nor g3380(n3395 ,n3384 ,n3390);
    xnor g3381(n3394 ,n4[3] ,n26[3]);
    nor g3382(n3676 ,n3384 ,n3382);
    xnor g3383(n3393 ,n4[2] ,n26[2]);
    xnor g3384(n3392 ,n4[5] ,n26[5]);
    xnor g3385(n3391 ,n4[4] ,n26[4]);
    xnor g3386(n3390 ,n4[1] ,n26[1]);
    xnor g3387(n3389 ,n4[6] ,n26[6]);
    xnor g3388(n3388 ,n4[7] ,n26[7]);
    nor g3389(n3387 ,n3371 ,n3375);
    nor g3390(n3386 ,n3372 ,n3369);
    nor g3391(n3385 ,n3370 ,n3378);
    nor g3392(n3384 ,n3373 ,n3374);
    nor g3393(n3383 ,n3376 ,n3377);
    nor g3394(n3382 ,n26[0] ,n4[0]);
    nor g3395(n3381 ,n26[6] ,n4[6]);
    nor g3396(n3380 ,n26[7] ,n4[7]);
    nor g3397(n3379 ,n26[1] ,n4[1]);
    not g3398(n3378 ,n4[4]);
    not g3399(n3377 ,n4[3]);
    not g3400(n3376 ,n26[3]);
    not g3401(n3375 ,n4[5]);
    not g3402(n3374 ,n4[0]);
    not g3403(n3373 ,n26[0]);
    not g3404(n3372 ,n26[2]);
    not g3405(n3371 ,n26[5]);
    not g3406(n3370 ,n26[4]);
    not g3407(n3369 ,n4[2]);
    xnor g3408(n3643 ,n3675 ,n3469);
    nor g3409(n3644 ,n3413 ,n3469);
    nor g3410(n3469 ,n3428 ,n3468);
    xnor g3411(n3642 ,n3442 ,n3466);
    nor g3412(n3468 ,n3442 ,n3467);
    not g3413(n3467 ,n3466);
    nor g3414(n3466 ,n3419 ,n3465);
    xnor g3415(n3641 ,n3437 ,n3464);
    nor g3416(n3465 ,n3437 ,n3464);
    nor g3417(n3464 ,n3422 ,n3463);
    xnor g3418(n3640 ,n3435 ,n3462);
    nor g3419(n3463 ,n3435 ,n3462);
    nor g3420(n3462 ,n3420 ,n3461);
    xnor g3421(n3685 ,n3432 ,n3460);
    nor g3422(n3461 ,n3432 ,n3460);
    nor g3423(n3460 ,n3425 ,n3459);
    xnor g3424(n3686 ,n3438 ,n3458);
    nor g3425(n3459 ,n3438 ,n3458);
    nor g3426(n3458 ,n3429 ,n3457);
    xnor g3427(n3687 ,n3431 ,n3456);
    nor g3428(n3457 ,n3431 ,n3456);
    nor g3429(n3456 ,n3426 ,n3455);
    xnor g3430(n3688 ,n3433 ,n3454);
    nor g3431(n3455 ,n3433 ,n3454);
    nor g3432(n3454 ,n3418 ,n3453);
    xnor g3433(n3689 ,n3434 ,n3452);
    nor g3434(n3453 ,n3434 ,n3452);
    nor g3435(n3452 ,n3421 ,n3451);
    xnor g3436(n3690 ,n3440 ,n3450);
    nor g3437(n3451 ,n3440 ,n3450);
    nor g3438(n3450 ,n3424 ,n3449);
    xor g3439(n3691 ,n3439 ,n3447);
    nor g3440(n3449 ,n3439 ,n3448);
    not g3441(n3448 ,n3447);
    nor g3442(n3447 ,n3427 ,n3446);
    xnor g3443(n3692 ,n3441 ,n3444);
    nor g3444(n3446 ,n3441 ,n3445);
    not g3445(n3445 ,n3444);
    nor g3446(n3444 ,n3417 ,n3443);
    xnor g3447(n3693 ,n3436 ,n3430);
    nor g3448(n3443 ,n3430 ,n3436);
    nor g3449(n3694 ,n3430 ,n3423);
    xnor g3450(n3442 ,n3674 ,n3661);
    xnor g3451(n3441 ,n3664 ,n3651);
    xnor g3452(n3440 ,n3666 ,n3653);
    xnor g3453(n3439 ,n3665 ,n3652);
    xnor g3454(n3438 ,n3670 ,n3657);
    xnor g3455(n3437 ,n3673 ,n3660);
    xnor g3456(n3436 ,n3650 ,n3663);
    xnor g3457(n3435 ,n3672 ,n3659);
    xnor g3458(n3434 ,n3667 ,n3654);
    xnor g3459(n3433 ,n3668 ,n3655);
    xnor g3460(n3432 ,n3671 ,n3658);
    xnor g3461(n3431 ,n3669 ,n3656);
    nor g3462(n3429 ,n3669 ,n3656);
    nor g3463(n3428 ,n3416 ,n3414);
    nor g3464(n3427 ,n3412 ,n3410);
    nor g3465(n3426 ,n3668 ,n3655);
    nor g3466(n3425 ,n3670 ,n3657);
    nor g3467(n3424 ,n3665 ,n3652);
    nor g3468(n3430 ,n3415 ,n3411);
    nor g3469(n3423 ,n3662 ,n3649);
    nor g3470(n3422 ,n3672 ,n3659);
    nor g3471(n3421 ,n3666 ,n3653);
    nor g3472(n3420 ,n3671 ,n3658);
    nor g3473(n3419 ,n3673 ,n3660);
    nor g3474(n3418 ,n3667 ,n3654);
    nor g3475(n3417 ,n3663 ,n3650);
    not g3476(n3416 ,n3674);
    not g3477(n3415 ,n3662);
    not g3478(n3414 ,n3661);
    not g3479(n3413 ,n3675);
    not g3480(n3412 ,n3664);
    not g3481(n3411 ,n3649);
    not g3482(n3410 ,n3651);
endmodule
