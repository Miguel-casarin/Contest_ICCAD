module top(n0, n1, n2, n3, n4, n5, n6);
    input n0, n1;
    input [13:0] n2;
    input [12:0] n3;
    output [12:0] n4, n5, n6;
    wire n0, n1;
    wire [13:0] n2;
    wire [12:0] n3;
    wire [12:0] n4, n5, n6;
    wire [12:0] n7;
    wire [12:0] n8;
    wire [12:0] n9;
    wire [12:0] n10;
    wire [12:0] n11;
    wire [12:0] n12;
    wire [12:0] n13;
    wire [2:0] n14;
    wire [3:0] n15;
    wire n16, n17, n18, n19, n20, n21, n22, n23;
    wire n24, n25, n26, n27, n28, n29, n30, n31;
    wire n32, n33, n34, n35, n36, n37, n38, n39;
    wire n40, n41, n42, n43, n44, n45, n46, n47;
    wire n48, n49, n50, n51, n52, n53, n54, n55;
    wire n56, n57, n58, n59, n60, n61, n62, n63;
    wire n64, n65, n66, n67, n68, n69, n70, n71;
    wire n72, n73, n74, n75, n76, n77, n78, n79;
    wire n80, n81, n82, n83, n84, n85, n86, n87;
    wire n88, n89, n90, n91, n92, n93, n94, n95;
    wire n96, n97, n98, n99, n100, n101, n102, n103;
    wire n104, n105, n106, n107, n108, n109, n110, n111;
    wire n112, n113, n114, n115, n116, n117, n118, n119;
    wire n120, n121, n122, n123, n124, n125, n126, n127;
    wire n128, n129, n130, n131, n132, n133, n134, n135;
    wire n136, n137, n138, n139, n140, n141, n142, n143;
    wire n144, n145, n146, n147, n148, n149, n150, n151;
    wire n152, n153, n154, n155, n156, n157, n158, n159;
    wire n160, n161, n162, n163, n164, n165, n166, n167;
    wire n168, n169, n170, n171, n172, n173, n174, n175;
    wire n176, n177, n178, n179, n180, n181, n182, n183;
    wire n184, n185, n186, n187, n188, n189, n190, n191;
    wire n192, n193, n194, n195, n196, n197, n198, n199;
    wire n200, n201, n202, n203, n204, n205, n206, n207;
    wire n208, n209, n210, n211, n212, n213, n214, n215;
    wire n216, n217, n218, n219, n220, n221, n222, n223;
    wire n224, n225, n226, n227, n228, n229, n230, n231;
    wire n232, n233, n234, n235, n236, n237, n238, n239;
    wire n240, n241, n242, n243, n244, n245, n246, n247;
    wire n248, n249, n250, n251, n252, n253, n254, n255;
    wire n256, n257, n258, n259, n260, n261, n262, n263;
    wire n264, n265, n266, n267, n268, n269, n270, n271;
    wire n272, n273, n274, n275, n276, n277, n278, n279;
    wire n280, n281, n282, n283, n284, n285, n286, n287;
    wire n288, n289, n290, n291, n292, n293, n294, n295;
    wire n296, n297, n298, n299, n300, n301, n302, n303;
    wire n304, n305, n306, n307, n308, n309, n310, n311;
    wire n312, n313, n314, n315, n316, n317, n318, n319;
    wire n320, n321, n322, n323, n324, n325, n326, n327;
    wire n328, n329, n330, n331, n332, n333, n334, n335;
    wire n336, n337, n338, n339, n340, n341, n342, n343;
    wire n344, n345, n346, n347, n348, n349, n350, n351;
    wire n352, n353, n354, n355, n356, n357, n358, n359;
    wire n360, n361, n362, n363, n364, n365, n366, n367;
    wire n368, n369, n370, n371, n372, n373, n374, n375;
    wire n376, n377, n378, n379, n380, n381, n382, n383;
    wire n384, n385, n386, n387, n388, n389, n390, n391;
    wire n392, n393, n394, n395, n396, n397, n398, n399;
    wire n400, n401, n402, n403, n404, n405, n406, n407;
    wire n408, n409, n410, n411, n412, n413, n414, n415;
    wire n416, n417, n418, n419, n420, n421, n422, n423;
    wire n424, n425, n426, n427, n428, n429, n430, n431;
    wire n432, n433, n434, n435, n436, n437, n438, n439;
    wire n440, n441, n442, n443, n444, n445, n446, n447;
    wire n448, n449, n450, n451, n452, n453, n454, n455;
    wire n456, n457, n458, n459, n460, n461, n462, n463;
    wire n464, n465, n466, n467, n468, n469, n470, n471;
    wire n472, n473, n474, n475, n476, n477, n478, n479;
    wire n480, n481, n482, n483, n484, n485, n486, n487;
    wire n488, n489, n490, n491, n492, n493, n494, n495;
    wire n496, n497, n498, n499, n500, n501, n502, n503;
    wire n504, n505, n506, n507, n508, n509, n510, n511;
    wire n512, n513, n514, n515, n516, n517, n518, n519;
    wire n520, n521, n522, n523, n524, n525, n526, n527;
    wire n528, n529, n530, n531, n532, n533, n534, n535;
    wire n536, n537, n538, n539, n540, n541, n542, n543;
    wire n544, n545, n546, n547, n548, n549, n550, n551;
    wire n552, n553, n554, n555, n556, n557, n558, n559;
    wire n560, n561, n562, n563, n564, n565, n566, n567;
    wire n568, n569, n570, n571, n572, n573, n574, n575;
    wire n576, n577, n578, n579, n580, n581, n582, n583;
    wire n584, n585, n586, n587, n588, n589, n590, n591;
    wire n592, n593, n594, n595, n596, n597, n598, n599;
    wire n600, n601, n602, n603, n604, n605, n606, n607;
    wire n608, n609, n610, n611, n612, n613, n614, n615;
    wire n616, n617, n618, n619, n620, n621, n622, n623;
    wire n624, n625, n626, n627, n628, n629, n630, n631;
    wire n632, n633, n634, n635, n636, n637, n638, n639;
    wire n640, n641, n642, n643, n644, n645, n646, n647;
    wire n648, n649, n650, n651, n652, n653, n654, n655;
    wire n656, n657, n658, n659, n660, n661, n662, n663;
    wire n664, n665, n666, n667, n668, n669, n670, n671;
    wire n672, n673, n674, n675, n676, n677, n678, n679;
    wire n680, n681, n682, n683, n684, n685, n686, n687;
    wire n688, n689, n690, n691, n692, n693, n694, n695;
    wire n696, n697, n698, n699, n700, n701, n702, n703;
    wire n704, n705, n706, n707, n708, n709, n710, n711;
    wire n712, n713, n714, n715, n716, n717, n718, n719;
    wire n720, n721, n722, n723, n724, n725, n726, n727;
    wire n728, n729, n730, n731, n732, n733, n734, n735;
    wire n736, n737, n738, n739, n740, n741, n742, n743;
    wire n744, n745, n746, n747, n748, n749, n750, n751;
    wire n752, n753, n754, n755, n756, n757, n758, n759;
    wire n760, n761, n762, n763, n764, n765, n766, n767;
    wire n768, n769, n770, n771, n772, n773, n774, n775;
    wire n776, n777, n778, n779, n780, n781, n782, n783;
    wire n784, n785, n786, n787, n788, n789, n790, n791;
    wire n792, n793, n794, n795, n796, n797, n798, n799;
    wire n800, n801, n802, n803, n804, n805, n806, n807;
    wire n808, n809, n810, n811, n812, n813, n814, n815;
    wire n816, n817, n818, n819, n820, n821, n822, n823;
    wire n824, n825, n826, n827, n828, n829, n830, n831;
    wire n832, n833, n834, n835, n836, n837, n838, n839;
    wire n840, n841, n842, n843, n844, n845, n846, n847;
    wire n848, n849;
    xnor g0(n5[3] ,n689 ,n8[3]);
    xnor g1(n4[10] ,n688 ,n9[10]);
    xnor g2(n4[9] ,n693 ,n9[9]);
    xnor g3(n4[6] ,n692 ,n9[6]);
    xnor g4(n4[5] ,n694 ,n9[5]);
    xnor g5(n5[11] ,n687 ,n8[11]);
    xnor g6(n5[10] ,n688 ,n8[10]);
    xnor g7(n5[9] ,n693 ,n8[9]);
    xnor g8(n5[8] ,n690 ,n8[8]);
    xnor g9(n4[8] ,n690 ,n9[8]);
    xnor g10(n5[7] ,n685 ,n8[7]);
    xnor g11(n5[6] ,n692 ,n8[6]);
    xnor g12(n5[5] ,n694 ,n8[5]);
    xnor g13(n5[4] ,n691 ,n8[4]);
    xnor g14(n4[4] ,n691 ,n9[4]);
    xnor g15(n4[11] ,n687 ,n9[11]);
    xnor g16(n5[2] ,n686 ,n8[2]);
    xnor g17(n5[1] ,n684 ,n8[1]);
    xnor g18(n4[7] ,n685 ,n9[7]);
    xnor g19(n4[3] ,n689 ,n9[3]);
    xnor g20(n6[11] ,n687 ,n10[11]);
    xnor g21(n6[10] ,n688 ,n10[10]);
    xnor g22(n6[9] ,n693 ,n10[9]);
    xnor g23(n4[2] ,n686 ,n9[2]);
    xnor g24(n6[8] ,n690 ,n10[8]);
    xnor g25(n6[7] ,n685 ,n10[7]);
    xnor g26(n6[6] ,n692 ,n10[6]);
    xnor g27(n6[5] ,n694 ,n10[5]);
    xnor g28(n4[1] ,n684 ,n9[1]);
    xnor g29(n6[4] ,n691 ,n10[4]);
    xnor g30(n6[3] ,n689 ,n10[3]);
    xnor g31(n6[2] ,n686 ,n10[2]);
    xnor g32(n6[1] ,n684 ,n10[1]);
    xnor g33(n4[0] ,n682 ,n9[0]);
    xnor g34(n5[12] ,n683 ,n8[12]);
    xnor g35(n5[0] ,n682 ,n8[0]);
    xnor g36(n6[12] ,n683 ,n10[12]);
    xnor g37(n4[12] ,n683 ,n9[12]);
    xnor g38(n6[0] ,n682 ,n10[0]);
    xnor g39(n694 ,n11[5] ,n680);
    xnor g40(n693 ,n11[9] ,n681);
    xnor g41(n692 ,n11[6] ,n671);
    xnor g42(n691 ,n11[4] ,n679);
    xnor g43(n690 ,n11[8] ,n678);
    xnor g44(n689 ,n11[3] ,n677);
    xnor g45(n688 ,n11[10] ,n676);
    xnor g46(n687 ,n11[11] ,n672);
    xnor g47(n686 ,n11[2] ,n675);
    xnor g48(n685 ,n11[7] ,n674);
    xnor g49(n684 ,n11[1] ,n673);
    xnor g50(n682 ,n3[0] ,n666);
    xor g51(n765 ,n11[9] ,n3[9]);
    xor g52(n764 ,n11[8] ,n3[8]);
    xor g53(n763 ,n11[7] ,n3[7]);
    xor g54(n762 ,n11[6] ,n3[6]);
    xor g55(n760 ,n11[4] ,n3[4]);
    xor g56(n759 ,n11[3] ,n3[3]);
    xor g57(n758 ,n11[2] ,n3[2]);
    xor g58(n757 ,n11[1] ,n3[1]);
    xor g59(n790 ,n11[8] ,n2[8]);
    xor g60(n789 ,n11[7] ,n2[7]);
    xor g61(n741 ,n11[11] ,n742);
    xor g62(n739 ,n11[10] ,n740);
    xor g63(n737 ,n11[9] ,n738);
    nor g64(n681 ,n702 ,n667);
    nor g65(n680 ,n706 ,n658);
    nor g66(n679 ,n701 ,n663);
    nor g67(n678 ,n704 ,n662);
    nor g68(n677 ,n695 ,n661);
    nor g69(n676 ,n705 ,n659);
    nor g70(n675 ,n703 ,n660);
    nor g71(n674 ,n699 ,n664);
    nor g72(n673 ,n700 ,n670);
    nor g73(n672 ,n707 ,n669);
    nor g74(n671 ,n696 ,n668);
    xor g75(n735 ,n11[8] ,n736);
    xor g76(n733 ,n11[7] ,n734);
    xor g77(n731 ,n11[6] ,n732);
    xor g78(n729 ,n11[5] ,n730);
    xor g79(n727 ,n11[4] ,n728);
    xor g80(n725 ,n11[3] ,n726);
    xor g81(n723 ,n11[2] ,n724);
    xor g82(n721 ,n11[1] ,n722);
    xor g83(n793 ,n11[11] ,n2[11]);
    xor g84(n792 ,n11[10] ,n2[10]);
    xor g85(n791 ,n11[9] ,n2[9]);
    xor g86(n784 ,n11[2] ,n2[2]);
    xor g87(n788 ,n11[6] ,n2[6]);
    xor g88(n786 ,n11[4] ,n2[4]);
    xor g89(n785 ,n11[3] ,n2[3]);
    xor g90(n783 ,n11[1] ,n2[1]);
    xor g91(n787 ,n11[5] ,n2[5]);
    xor g92(n761 ,n11[5] ,n3[5]);
    xor g93(n767 ,n11[11] ,n3[11]);
    xor g94(n766 ,n11[10] ,n3[10]);
    xor g95(n782 ,n2[0] ,n3[0]);
    not g96(n13[1] ,n670);
    not g97(n13[11] ,n669);
    not g98(n13[6] ,n668);
    not g99(n13[9] ,n667);
    nor g100(n666 ,n657 ,n698);
    nor g101(n665 ,n656 ,n697);
    nor g102(n670 ,n3[0] ,n11[2]);
    nor g103(n668 ,n11[7] ,n11[5]);
    nor g104(n667 ,n11[10] ,n11[8]);
    not g105(n13[7] ,n664);
    not g106(n13[4] ,n663);
    not g107(n13[8] ,n662);
    not g108(n13[3] ,n661);
    not g109(n13[2] ,n660);
    not g110(n13[10] ,n659);
    not g111(n13[5] ,n658);
    nor g112(n664 ,n11[8] ,n11[6]);
    nor g113(n663 ,n11[5] ,n11[3]);
    nor g114(n662 ,n11[9] ,n11[7]);
    nor g115(n661 ,n11[4] ,n11[2]);
    nor g116(n660 ,n11[3] ,n11[1]);
    nor g117(n659 ,n11[11] ,n11[9]);
    nor g118(n658 ,n11[6] ,n11[4]);
    not g119(n657 ,n11[1]);
    not g120(n656 ,n11[11]);
    dff g121(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n595), .Q(n9[0]));
    dff g122(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n571), .Q(n9[1]));
    dff g123(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n604), .Q(n9[2]));
    dff g124(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n598), .Q(n9[3]));
    dff g125(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n597), .Q(n9[4]));
    dff g126(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n588), .Q(n9[5]));
    dff g127(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n587), .Q(n9[6]));
    dff g128(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n582), .Q(n9[7]));
    dff g129(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n581), .Q(n9[8]));
    dff g130(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n580), .Q(n9[9]));
    dff g131(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n576), .Q(n9[10]));
    dff g132(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n579), .Q(n9[11]));
    dff g133(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n578), .Q(n9[12]));
    dff g134(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n577), .Q(n8[0]));
    dff g135(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n602), .Q(n8[1]));
    dff g136(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n575), .Q(n8[2]));
    dff g137(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n574), .Q(n8[3]));
    dff g138(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n573), .Q(n8[4]));
    dff g139(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n572), .Q(n8[5]));
    dff g140(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n603), .Q(n8[6]));
    dff g141(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n617), .Q(n8[7]));
    dff g142(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n632), .Q(n8[8]));
    dff g143(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n568), .Q(n8[9]));
    dff g144(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n601), .Q(n8[10]));
    dff g145(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n600), .Q(n8[11]));
    dff g146(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n599), .Q(n8[12]));
    dff g147(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n641), .Q(n10[0]));
    dff g148(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n569), .Q(n10[1]));
    dff g149(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n596), .Q(n10[2]));
    dff g150(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n594), .Q(n10[3]));
    dff g151(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n593), .Q(n10[4]));
    dff g152(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n592), .Q(n10[5]));
    dff g153(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n591), .Q(n10[6]));
    dff g154(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n590), .Q(n10[7]));
    dff g155(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n589), .Q(n10[8]));
    dff g156(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n586), .Q(n10[9]));
    dff g157(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n585), .Q(n10[10]));
    dff g158(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n584), .Q(n10[11]));
    dff g159(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n583), .Q(n10[12]));
    dff g160(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n497), .Q(n14[0]));
    dff g161(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n496), .Q(n14[1]));
    dff g162(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n526), .Q(n14[2]));
    dff g163(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n655), .Q(n15[0]));
    dff g164(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n654), .Q(n15[1]));
    dff g165(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n653), .Q(n15[2]));
    nor g166(n655 ,n1 ,n652);
    nor g167(n654 ,n1 ,n651);
    nor g168(n653 ,n1 ,n649);
    or g169(n652 ,n365 ,n650);
    or g170(n651 ,n374 ,n650);
    not g171(n649 ,n650);
    nor g172(n650 ,n370 ,n634);
    or g173(n648 ,n619 ,n618);
    or g174(n647 ,n630 ,n629);
    or g175(n646 ,n627 ,n628);
    or g176(n645 ,n626 ,n625);
    or g177(n644 ,n623 ,n624);
    or g178(n643 ,n620 ,n622);
    or g179(n642 ,n631 ,n621);
    or g180(n641 ,n558 ,n570);
    or g181(n640 ,n616 ,n633);
    or g182(n639 ,n615 ,n614);
    or g183(n638 ,n612 ,n613);
    or g184(n637 ,n611 ,n610);
    or g185(n636 ,n608 ,n609);
    or g186(n635 ,n606 ,n607);
    nor g187(n634 ,n15[0] ,n605);
    nor g188(n633 ,n260 ,n567);
    or g189(n632 ,n564 ,n524);
    nor g190(n631 ,n308 ,n527);
    nor g191(n630 ,n318 ,n527);
    nor g192(n629 ,n252 ,n567);
    nor g193(n628 ,n263 ,n567);
    nor g194(n627 ,n314 ,n527);
    nor g195(n626 ,n320 ,n527);
    nor g196(n625 ,n258 ,n567);
    nor g197(n624 ,n255 ,n567);
    nor g198(n623 ,n313 ,n527);
    nor g199(n622 ,n256 ,n567);
    nor g200(n621 ,n265 ,n567);
    nor g201(n620 ,n316 ,n527);
    nor g202(n619 ,n310 ,n527);
    nor g203(n618 ,n253 ,n567);
    or g204(n617 ,n565 ,n525);
    nor g205(n616 ,n319 ,n527);
    nor g206(n615 ,n311 ,n527);
    nor g207(n614 ,n261 ,n567);
    nor g208(n613 ,n259 ,n567);
    nor g209(n612 ,n312 ,n527);
    nor g210(n611 ,n317 ,n527);
    nor g211(n610 ,n254 ,n567);
    nor g212(n609 ,n262 ,n567);
    nor g213(n608 ,n315 ,n527);
    nor g214(n607 ,n266 ,n567);
    nor g215(n606 ,n307 ,n527);
    nor g216(n605 ,n361 ,n530);
    or g217(n604 ,n561 ,n518);
    or g218(n603 ,n546 ,n528);
    or g219(n602 ,n428 ,n490);
    or g220(n601 ,n562 ,n520);
    or g221(n600 ,n560 ,n519);
    or g222(n599 ,n559 ,n517);
    or g223(n598 ,n557 ,n516);
    or g224(n597 ,n554 ,n512);
    or g225(n596 ,n556 ,n514);
    or g226(n595 ,n539 ,n492);
    or g227(n594 ,n555 ,n513);
    or g228(n593 ,n553 ,n491);
    or g229(n592 ,n552 ,n511);
    or g230(n591 ,n550 ,n510);
    or g231(n590 ,n549 ,n508);
    or g232(n589 ,n548 ,n507);
    or g233(n588 ,n551 ,n509);
    or g234(n587 ,n566 ,n505);
    or g235(n586 ,n547 ,n506);
    or g236(n585 ,n545 ,n523);
    or g237(n584 ,n544 ,n504);
    or g238(n583 ,n543 ,n503);
    or g239(n582 ,n542 ,n501);
    or g240(n581 ,n541 ,n499);
    or g241(n580 ,n540 ,n498);
    or g242(n579 ,n537 ,n495);
    or g243(n578 ,n536 ,n494);
    or g244(n577 ,n535 ,n493);
    or g245(n576 ,n538 ,n500);
    or g246(n575 ,n534 ,n489);
    or g247(n574 ,n533 ,n488);
    or g248(n573 ,n532 ,n487);
    or g249(n572 ,n531 ,n502);
    or g250(n571 ,n460 ,n522);
    or g251(n570 ,n480 ,n529);
    or g252(n569 ,n453 ,n515);
    or g253(n568 ,n563 ,n521);
    nor g254(n566 ,n324 ,n436);
    nor g255(n565 ,n358 ,n448);
    nor g256(n564 ,n353 ,n447);
    nor g257(n563 ,n357 ,n443);
    nor g258(n562 ,n334 ,n444);
    nor g259(n561 ,n344 ,n441);
    nor g260(n560 ,n264 ,n442);
    nor g261(n559 ,n332 ,n440);
    nor g262(n558 ,n347 ,n437);
    nor g263(n557 ,n342 ,n439);
    nor g264(n556 ,n341 ,n441);
    nor g265(n555 ,n333 ,n439);
    nor g266(n554 ,n336 ,n445);
    nor g267(n553 ,n350 ,n445);
    nor g268(n552 ,n325 ,n446);
    nor g269(n551 ,n345 ,n446);
    nor g270(n550 ,n328 ,n436);
    nor g271(n549 ,n331 ,n448);
    nor g272(n548 ,n339 ,n447);
    nor g273(n547 ,n349 ,n443);
    nor g274(n546 ,n326 ,n436);
    nor g275(n545 ,n327 ,n444);
    nor g276(n544 ,n354 ,n442);
    nor g277(n543 ,n351 ,n440);
    nor g278(n542 ,n330 ,n448);
    nor g279(n541 ,n335 ,n447);
    nor g280(n540 ,n356 ,n443);
    nor g281(n539 ,n348 ,n437);
    nor g282(n538 ,n337 ,n444);
    nor g283(n537 ,n343 ,n442);
    nor g284(n536 ,n329 ,n440);
    nor g285(n535 ,n340 ,n437);
    nor g286(n534 ,n352 ,n441);
    nor g287(n533 ,n355 ,n439);
    nor g288(n532 ,n346 ,n445);
    nor g289(n531 ,n338 ,n446);
    or g290(n530 ,n378 ,n421);
    nor g291(n529 ,n368 ,n420);
    or g292(n528 ,n462 ,n479);
    or g293(n567 ,n1 ,n450);
    nor g294(n526 ,n1 ,n416);
    or g295(n525 ,n461 ,n486);
    or g296(n524 ,n459 ,n481);
    or g297(n523 ,n474 ,n483);
    nor g298(n522 ,n419 ,n438);
    or g299(n521 ,n468 ,n482);
    or g300(n520 ,n457 ,n483);
    or g301(n519 ,n431 ,n484);
    or g302(n518 ,n454 ,n475);
    or g303(n517 ,n455 ,n485);
    or g304(n516 ,n451 ,n477);
    nor g305(n515 ,n417 ,n438);
    or g306(n514 ,n458 ,n475);
    or g307(n513 ,n456 ,n477);
    or g308(n512 ,n465 ,n478);
    or g309(n511 ,n466 ,n476);
    or g310(n510 ,n467 ,n479);
    or g311(n509 ,n463 ,n476);
    or g312(n508 ,n470 ,n486);
    or g313(n507 ,n469 ,n481);
    or g314(n506 ,n452 ,n482);
    or g315(n505 ,n472 ,n479);
    or g316(n504 ,n471 ,n484);
    or g317(n503 ,n473 ,n485);
    or g318(n502 ,n423 ,n476);
    or g319(n501 ,n418 ,n486);
    or g320(n500 ,n434 ,n483);
    or g321(n499 ,n422 ,n481);
    or g322(n498 ,n433 ,n482);
    nor g323(n497 ,n1 ,n435);
    nor g324(n496 ,n1 ,n414);
    or g325(n495 ,n432 ,n484);
    or g326(n494 ,n430 ,n485);
    or g327(n493 ,n429 ,n480);
    or g328(n492 ,n427 ,n480);
    or g329(n491 ,n464 ,n478);
    nor g330(n490 ,n415 ,n438);
    or g331(n489 ,n426 ,n475);
    or g332(n488 ,n425 ,n477);
    or g333(n487 ,n424 ,n478);
    or g334(n527 ,n1 ,n449);
    nor g335(n474 ,n290 ,n385);
    nor g336(n473 ,n273 ,n385);
    nor g337(n472 ,n276 ,n385);
    nor g338(n471 ,n272 ,n385);
    nor g339(n470 ,n306 ,n385);
    nor g340(n469 ,n288 ,n385);
    nor g341(n468 ,n298 ,n385);
    nor g342(n467 ,n289 ,n385);
    nor g343(n466 ,n294 ,n385);
    nor g344(n465 ,n303 ,n385);
    nor g345(n464 ,n267 ,n385);
    nor g346(n463 ,n280 ,n385);
    nor g347(n462 ,n302 ,n385);
    nor g348(n461 ,n284 ,n385);
    nor g349(n460 ,n278 ,n385);
    nor g350(n459 ,n281 ,n385);
    nor g351(n458 ,n274 ,n385);
    nor g352(n457 ,n286 ,n385);
    nor g353(n456 ,n285 ,n385);
    nor g354(n455 ,n304 ,n385);
    nor g355(n454 ,n301 ,n385);
    nor g356(n453 ,n271 ,n385);
    nor g357(n452 ,n300 ,n385);
    nor g358(n451 ,n269 ,n385);
    nor g359(n486 ,n319 ,n409);
    nor g360(n485 ,n307 ,n395);
    nor g361(n484 ,n315 ,n407);
    nor g362(n483 ,n317 ,n405);
    nor g363(n482 ,n312 ,n397);
    nor g364(n481 ,n311 ,n391);
    nor g365(n480 ,n318 ,n389);
    nor g366(n479 ,n310 ,n393);
    nor g367(n478 ,n316 ,n387);
    nor g368(n477 ,n313 ,n413);
    nor g369(n476 ,n308 ,n411);
    nor g370(n475 ,n320 ,n403);
    not g371(n450 ,n449);
    xnor g372(n435 ,n377 ,n14[0]);
    nor g373(n434 ,n305 ,n385);
    nor g374(n433 ,n277 ,n385);
    nor g375(n432 ,n275 ,n385);
    nor g376(n431 ,n279 ,n385);
    nor g377(n430 ,n296 ,n385);
    nor g378(n429 ,n291 ,n385);
    nor g379(n428 ,n283 ,n385);
    nor g380(n427 ,n270 ,n385);
    nor g381(n426 ,n268 ,n385);
    nor g382(n425 ,n282 ,n385);
    nor g383(n424 ,n292 ,n385);
    nor g384(n423 ,n293 ,n385);
    nor g385(n422 ,n299 ,n385);
    or g386(n421 ,n366 ,n384);
    or g387(n420 ,n363 ,n385);
    nor g388(n419 ,n9[1] ,n401);
    nor g389(n418 ,n287 ,n385);
    nor g390(n417 ,n10[1] ,n401);
    nor g391(n416 ,n382 ,n399);
    nor g392(n415 ,n8[1] ,n401);
    nor g393(n414 ,n383 ,n400);
    nor g394(n449 ,n362 ,n381);
    nor g395(n448 ,n375 ,n408);
    nor g396(n447 ,n375 ,n390);
    nor g397(n446 ,n375 ,n410);
    nor g398(n445 ,n375 ,n386);
    nor g399(n444 ,n375 ,n404);
    nor g400(n443 ,n375 ,n396);
    nor g401(n442 ,n375 ,n406);
    nor g402(n441 ,n375 ,n402);
    nor g403(n440 ,n375 ,n394);
    nor g404(n439 ,n375 ,n412);
    nor g405(n438 ,n375 ,n398);
    nor g406(n437 ,n375 ,n388);
    nor g407(n436 ,n375 ,n392);
    not g408(n413 ,n412);
    not g409(n411 ,n410);
    not g410(n409 ,n408);
    not g411(n407 ,n406);
    not g412(n405 ,n404);
    not g413(n403 ,n402);
    nor g414(n400 ,n297 ,n376);
    nor g415(n399 ,n295 ,n376);
    nor g416(n398 ,n263 ,n380);
    nor g417(n412 ,n255 ,n380);
    nor g418(n410 ,n265 ,n380);
    nor g419(n408 ,n260 ,n380);
    nor g420(n406 ,n262 ,n380);
    nor g421(n404 ,n254 ,n380);
    nor g422(n402 ,n258 ,n380);
    nor g423(n401 ,n314 ,n380);
    not g424(n397 ,n396);
    not g425(n395 ,n394);
    not g426(n393 ,n392);
    not g427(n391 ,n390);
    not g428(n389 ,n388);
    not g429(n387 ,n386);
    nor g430(n383 ,n321 ,n377);
    nor g431(n382 ,n322 ,n377);
    or g432(n381 ,n14[2] ,n376);
    nor g433(n396 ,n259 ,n380);
    nor g434(n394 ,n266 ,n380);
    nor g435(n392 ,n253 ,n380);
    nor g436(n390 ,n261 ,n380);
    nor g437(n388 ,n252 ,n380);
    nor g438(n386 ,n256 ,n380);
    or g439(n385 ,n15[2] ,n373);
    or g440(n379 ,n367 ,n360);
    or g441(n378 ,n359 ,n364);
    or g442(n380 ,n370 ,n371);
    not g443(n376 ,n377);
    nor g444(n374 ,n372 ,n369);
    or g445(n373 ,n15[1] ,n371);
    nor g446(n377 ,n15[1] ,n365);
    nor g447(n375 ,n1 ,n372);
    not g448(n370 ,n369);
    nor g449(n368 ,n252 ,n257);
    nor g450(n372 ,n309 ,n15[2]);
    or g451(n371 ,n309 ,n1);
    nor g452(n369 ,n323 ,n15[2]);
    nor g453(n363 ,n3[0] ,n708);
    or g454(n362 ,n14[0] ,n14[1]);
    or g455(n365 ,n15[0] ,n15[2]);
    not g456(n358 ,n8[7]);
    not g457(n357 ,n8[9]);
    not g458(n356 ,n9[9]);
    not g459(n355 ,n8[3]);
    not g460(n354 ,n10[11]);
    not g461(n353 ,n8[8]);
    not g462(n352 ,n8[2]);
    not g463(n351 ,n10[12]);
    not g464(n350 ,n10[4]);
    not g465(n349 ,n10[9]);
    not g466(n348 ,n9[0]);
    not g467(n347 ,n10[0]);
    not g468(n346 ,n8[4]);
    not g469(n345 ,n9[5]);
    not g470(n344 ,n9[2]);
    not g471(n343 ,n9[11]);
    not g472(n342 ,n9[3]);
    not g473(n341 ,n10[2]);
    not g474(n340 ,n8[0]);
    not g475(n339 ,n10[8]);
    not g476(n338 ,n8[5]);
    not g477(n337 ,n9[10]);
    not g478(n336 ,n9[4]);
    not g479(n335 ,n9[8]);
    not g480(n334 ,n8[10]);
    not g481(n333 ,n10[3]);
    not g482(n332 ,n8[12]);
    not g483(n331 ,n10[7]);
    not g484(n330 ,n9[7]);
    not g485(n329 ,n9[12]);
    not g486(n328 ,n10[6]);
    not g487(n327 ,n10[10]);
    not g488(n326 ,n8[6]);
    not g489(n325 ,n10[5]);
    not g490(n324 ,n9[6]);
    not g491(n323 ,n15[1]);
    not g492(n322 ,n14[2]);
    not g493(n321 ,n14[1]);
    not g494(n309 ,n15[0]);
    not g495(n306 ,n715);
    not g496(n305 ,n779);
    not g497(n304 ,n756);
    not g498(n303 ,n773);
    not g499(n302 ,n750);
    not g500(n301 ,n771);
    not g501(n300 ,n717);
    not g502(n299 ,n777);
    not g503(n298 ,n753);
    not g504(n297 ,n796);
    not g505(n296 ,n781);
    not g506(n295 ,n795);
    not g507(n294 ,n713);
    not g508(n293 ,n749);
    not g509(n292 ,n748);
    not g510(n291 ,n13[1]);
    not g511(n290 ,n718);
    not g512(n289 ,n714);
    not g513(n288 ,n716);
    not g514(n287 ,n776);
    not g515(n286 ,n754);
    not g516(n285 ,n711);
    not g517(n284 ,n751);
    not g518(n283 ,n745);
    not g519(n282 ,n747);
    not g520(n281 ,n752);
    not g521(n280 ,n774);
    not g522(n279 ,n755);
    not g523(n278 ,n770);
    not g524(n277 ,n778);
    not g525(n276 ,n775);
    not g526(n275 ,n780);
    not g527(n274 ,n710);
    not g528(n273 ,n720);
    not g529(n272 ,n719);
    not g530(n271 ,n709);
    not g531(n270 ,n769);
    not g532(n269 ,n772);
    not g533(n268 ,n746);
    not g534(n267 ,n712);
    not g535(n265 ,n11[5]);
    not g536(n264 ,n8[11]);
    not g537(n263 ,n11[1]);
    not g538(n262 ,n11[11]);
    not g539(n261 ,n11[8]);
    not g540(n260 ,n11[7]);
    not g541(n259 ,n11[9]);
    not g542(n258 ,n11[2]);
    not g543(n257 ,n708);
    not g544(n256 ,n11[4]);
    not g545(n255 ,n11[3]);
    not g546(n254 ,n11[10]);
    not g547(n253 ,n11[6]);
    not g548(n252 ,n3[0]);
    xnor g549(n781 ,n794 ,n82);
    nor g550(n82 ,n43 ,n81);
    xor g551(n780 ,n57 ,n80);
    nor g552(n81 ,n57 ,n80);
    nor g553(n80 ,n40 ,n79);
    xor g554(n779 ,n55 ,n78);
    nor g555(n79 ,n55 ,n78);
    nor g556(n78 ,n46 ,n77);
    xor g557(n778 ,n53 ,n76);
    nor g558(n77 ,n53 ,n76);
    nor g559(n76 ,n36 ,n75);
    xor g560(n777 ,n51 ,n74);
    nor g561(n75 ,n51 ,n74);
    nor g562(n74 ,n47 ,n73);
    xor g563(n776 ,n56 ,n72);
    nor g564(n73 ,n56 ,n72);
    nor g565(n72 ,n45 ,n71);
    xor g566(n775 ,n54 ,n70);
    nor g567(n71 ,n54 ,n70);
    nor g568(n70 ,n44 ,n69);
    xor g569(n774 ,n58 ,n68);
    nor g570(n69 ,n58 ,n68);
    nor g571(n68 ,n41 ,n67);
    xor g572(n773 ,n52 ,n66);
    nor g573(n67 ,n52 ,n66);
    nor g574(n66 ,n39 ,n65);
    xnor g575(n772 ,n59 ,n63);
    nor g576(n65 ,n59 ,n64);
    not g577(n64 ,n63);
    nor g578(n63 ,n38 ,n62);
    xnor g579(n771 ,n50 ,n61);
    nor g580(n62 ,n50 ,n61);
    nor g581(n61 ,n37 ,n60);
    xnor g582(n770 ,n49 ,n48);
    nor g583(n60 ,n48 ,n49);
    nor g584(n769 ,n48 ,n42);
    xnor g585(n59 ,n785 ,n13[3]);
    xnor g586(n58 ,n787 ,n13[5]);
    xnor g587(n57 ,n793 ,n13[11]);
    xnor g588(n56 ,n789 ,n13[7]);
    xnor g589(n55 ,n792 ,n13[10]);
    xnor g590(n54 ,n788 ,n13[6]);
    xnor g591(n53 ,n791 ,n13[9]);
    xnor g592(n52 ,n786 ,n13[4]);
    xnor g593(n51 ,n790 ,n13[8]);
    xnor g594(n50 ,n784 ,n13[2]);
    xnor g595(n49 ,n783 ,n13[1]);
    nor g596(n47 ,n17 ,n25);
    nor g597(n46 ,n33 ,n34);
    nor g598(n45 ,n30 ,n29);
    nor g599(n44 ,n31 ,n21);
    nor g600(n43 ,n28 ,n20);
    nor g601(n48 ,n18 ,n16);
    nor g602(n42 ,n782 ,n11[1]);
    nor g603(n41 ,n19 ,n26);
    nor g604(n40 ,n32 ,n35);
    nor g605(n39 ,n22 ,n23);
    nor g606(n38 ,n784 ,n13[2]);
    nor g607(n37 ,n783 ,n13[1]);
    nor g608(n36 ,n24 ,n27);
    not g609(n35 ,n13[10]);
    not g610(n34 ,n13[9]);
    not g611(n33 ,n791);
    not g612(n32 ,n792);
    not g613(n31 ,n787);
    not g614(n30 ,n788);
    not g615(n29 ,n13[6]);
    not g616(n28 ,n793);
    not g617(n27 ,n13[8]);
    not g618(n26 ,n13[4]);
    not g619(n25 ,n13[7]);
    not g620(n24 ,n790);
    not g621(n23 ,n13[3]);
    not g622(n22 ,n785);
    not g623(n21 ,n13[5]);
    not g624(n20 ,n13[11]);
    not g625(n19 ,n786);
    not g626(n18 ,n782);
    not g627(n17 ,n789);
    not g628(n16 ,n11[1]);
    xor g629(n756 ,n768 ,n130);
    nor g630(n130 ,n94 ,n129);
    xnor g631(n755 ,n106 ,n128);
    nor g632(n129 ,n106 ,n128);
    nor g633(n128 ,n88 ,n127);
    xor g634(n754 ,n108 ,n125);
    nor g635(n127 ,n108 ,n126);
    not g636(n126 ,n125);
    nor g637(n125 ,n95 ,n124);
    xnor g638(n753 ,n107 ,n122);
    nor g639(n124 ,n107 ,n123);
    not g640(n123 ,n122);
    nor g641(n122 ,n90 ,n121);
    xnor g642(n752 ,n99 ,n120);
    nor g643(n121 ,n99 ,n120);
    nor g644(n120 ,n92 ,n119);
    xnor g645(n751 ,n105 ,n118);
    nor g646(n119 ,n105 ,n118);
    nor g647(n118 ,n93 ,n117);
    xnor g648(n750 ,n102 ,n116);
    nor g649(n117 ,n102 ,n116);
    nor g650(n116 ,n91 ,n115);
    xnor g651(n749 ,n101 ,n114);
    nor g652(n115 ,n101 ,n114);
    nor g653(n114 ,n89 ,n113);
    xnor g654(n748 ,n100 ,n112);
    nor g655(n113 ,n100 ,n112);
    nor g656(n112 ,n87 ,n111);
    xnor g657(n747 ,n103 ,n110);
    nor g658(n111 ,n103 ,n110);
    nor g659(n110 ,n96 ,n109);
    xnor g660(n746 ,n104 ,n98);
    nor g661(n109 ,n98 ,n104);
    nor g662(n745 ,n98 ,n97);
    xnor g663(n108 ,n766 ,n13[11]);
    xnor g664(n107 ,n765 ,n13[10]);
    xnor g665(n106 ,n767 ,n11[11]);
    xnor g666(n105 ,n763 ,n13[8]);
    xnor g667(n104 ,n758 ,n13[3]);
    xnor g668(n103 ,n759 ,n13[4]);
    xnor g669(n102 ,n762 ,n13[7]);
    xnor g670(n101 ,n761 ,n13[6]);
    xnor g671(n100 ,n760 ,n13[5]);
    xnor g672(n99 ,n764 ,n13[9]);
    nor g673(n97 ,n757 ,n13[2]);
    nor g674(n96 ,n758 ,n13[3]);
    nor g675(n95 ,n84 ,n86);
    nor g676(n94 ,n767 ,n11[11]);
    nor g677(n93 ,n762 ,n13[7]);
    nor g678(n98 ,n83 ,n85);
    nor g679(n92 ,n763 ,n13[8]);
    nor g680(n91 ,n761 ,n13[6]);
    nor g681(n90 ,n764 ,n13[9]);
    nor g682(n89 ,n760 ,n13[5]);
    nor g683(n88 ,n766 ,n13[11]);
    nor g684(n87 ,n759 ,n13[4]);
    not g685(n86 ,n13[10]);
    not g686(n85 ,n13[2]);
    not g687(n84 ,n765);
    not g688(n83 ,n757);
    xnor g689(n744 ,n150 ,n185);
    nor g690(n185 ,n138 ,n184);
    xnor g691(n742 ,n156 ,n183);
    nor g692(n184 ,n156 ,n183);
    nor g693(n183 ,n144 ,n182);
    xnor g694(n740 ,n154 ,n181);
    nor g695(n182 ,n154 ,n181);
    nor g696(n181 ,n139 ,n180);
    xnor g697(n738 ,n153 ,n179);
    nor g698(n180 ,n153 ,n179);
    nor g699(n179 ,n141 ,n178);
    xor g700(n736 ,n159 ,n176);
    nor g701(n178 ,n159 ,n177);
    not g702(n177 ,n176);
    nor g703(n176 ,n148 ,n175);
    xor g704(n734 ,n160 ,n174);
    nor g705(n175 ,n160 ,n174);
    nor g706(n174 ,n146 ,n173);
    xnor g707(n732 ,n161 ,n171);
    nor g708(n173 ,n161 ,n172);
    not g709(n172 ,n171);
    nor g710(n171 ,n140 ,n170);
    xnor g711(n730 ,n155 ,n169);
    nor g712(n170 ,n155 ,n169);
    nor g713(n169 ,n142 ,n168);
    xnor g714(n728 ,n152 ,n167);
    nor g715(n168 ,n152 ,n167);
    nor g716(n167 ,n145 ,n166);
    xnor g717(n726 ,n158 ,n165);
    nor g718(n166 ,n158 ,n165);
    nor g719(n165 ,n137 ,n164);
    xnor g720(n724 ,n157 ,n163);
    nor g721(n164 ,n157 ,n163);
    nor g722(n163 ,n147 ,n162);
    xnor g723(n722 ,n151 ,n149);
    nor g724(n162 ,n149 ,n151);
    nor g725(n708 ,n149 ,n143);
    xnor g726(n161 ,n2[6] ,n3[6]);
    xnor g727(n160 ,n2[7] ,n3[7]);
    xnor g728(n159 ,n2[8] ,n3[8]);
    xnor g729(n158 ,n2[3] ,n3[3]);
    xnor g730(n157 ,n2[2] ,n3[2]);
    xnor g731(n150 ,n2[12] ,n3[12]);
    xnor g732(n156 ,n2[11] ,n3[11]);
    xnor g733(n155 ,n2[5] ,n3[5]);
    xnor g734(n154 ,n2[10] ,n3[10]);
    xnor g735(n153 ,n2[9] ,n3[9]);
    xnor g736(n152 ,n2[4] ,n3[4]);
    xnor g737(n151 ,n2[1] ,n3[1]);
    nor g738(n148 ,n135 ,n136);
    nor g739(n147 ,n2[1] ,n3[1]);
    nor g740(n146 ,n133 ,n132);
    nor g741(n145 ,n2[3] ,n3[3]);
    nor g742(n144 ,n2[10] ,n3[10]);
    nor g743(n149 ,n134 ,n131);
    nor g744(n143 ,n2[0] ,n3[0]);
    nor g745(n142 ,n2[4] ,n3[4]);
    nor g746(n141 ,n2[8] ,n3[8]);
    nor g747(n140 ,n2[5] ,n3[5]);
    nor g748(n139 ,n2[9] ,n3[9]);
    nor g749(n138 ,n2[11] ,n3[11]);
    nor g750(n137 ,n2[2] ,n3[2]);
    not g751(n136 ,n3[7]);
    not g752(n135 ,n2[7]);
    not g753(n134 ,n2[0]);
    not g754(n133 ,n2[6]);
    not g755(n132 ,n3[6]);
    not g756(n131 ,n3[0]);
    xor g757(n720 ,n216 ,n247);
    nor g758(n247 ,n211 ,n246);
    xor g759(n719 ,n222 ,n245);
    nor g760(n246 ,n222 ,n245);
    nor g761(n245 ,n214 ,n244);
    xor g762(n718 ,n224 ,n243);
    nor g763(n244 ,n224 ,n243);
    nor g764(n243 ,n210 ,n242);
    xor g765(n717 ,n221 ,n241);
    nor g766(n242 ,n221 ,n241);
    nor g767(n241 ,n207 ,n240);
    xor g768(n716 ,n223 ,n239);
    nor g769(n240 ,n223 ,n239);
    nor g770(n239 ,n213 ,n238);
    xor g771(n715 ,n226 ,n237);
    nor g772(n238 ,n226 ,n237);
    nor g773(n237 ,n204 ,n236);
    xor g774(n714 ,n225 ,n235);
    nor g775(n236 ,n225 ,n235);
    nor g776(n235 ,n212 ,n234);
    xor g777(n713 ,n220 ,n233);
    nor g778(n234 ,n220 ,n233);
    nor g779(n233 ,n208 ,n232);
    xnor g780(n712 ,n219 ,n230);
    nor g781(n232 ,n219 ,n231);
    not g782(n231 ,n230);
    nor g783(n230 ,n206 ,n229);
    xnor g784(n711 ,n218 ,n228);
    nor g785(n229 ,n218 ,n228);
    nor g786(n228 ,n205 ,n227);
    xnor g787(n710 ,n217 ,n215);
    nor g788(n227 ,n215 ,n217);
    nor g789(n709 ,n215 ,n209);
    xnor g790(n226 ,n733 ,n13[6]);
    xnor g791(n225 ,n731 ,n13[5]);
    xnor g792(n224 ,n739 ,n13[9]);
    xnor g793(n223 ,n735 ,n13[7]);
    xnor g794(n222 ,n741 ,n13[10]);
    xnor g795(n221 ,n737 ,n13[8]);
    xnor g796(n220 ,n729 ,n13[4]);
    xnor g797(n219 ,n727 ,n13[3]);
    xnor g798(n218 ,n725 ,n13[2]);
    xnor g799(n217 ,n723 ,n13[1]);
    xnor g800(n216 ,n13[11] ,n743);
    nor g801(n214 ,n202 ,n187);
    nor g802(n213 ,n199 ,n195);
    nor g803(n212 ,n188 ,n189);
    nor g804(n211 ,n200 ,n186);
    nor g805(n210 ,n201 ,n203);
    nor g806(n215 ,n192 ,n190);
    nor g807(n209 ,n721 ,n11[1]);
    nor g808(n208 ,n191 ,n198);
    nor g809(n207 ,n196 ,n194);
    nor g810(n206 ,n725 ,n13[2]);
    nor g811(n205 ,n723 ,n13[1]);
    nor g812(n204 ,n193 ,n197);
    not g813(n203 ,n13[8]);
    not g814(n202 ,n739);
    not g815(n201 ,n737);
    not g816(n200 ,n741);
    not g817(n199 ,n733);
    not g818(n198 ,n13[3]);
    not g819(n197 ,n13[5]);
    not g820(n196 ,n735);
    not g821(n195 ,n13[6]);
    not g822(n194 ,n13[7]);
    not g823(n193 ,n731);
    not g824(n192 ,n721);
    not g825(n191 ,n727);
    not g826(n190 ,n11[1]);
    not g827(n189 ,n13[4]);
    not g828(n188 ,n729);
    not g829(n187 ,n13[9]);
    not g830(n186 ,n13[10]);
    xor g831(n795 ,n14[2] ,n251);
    nor g832(n796 ,n251 ,n250);
    nor g833(n251 ,n249 ,n248);
    nor g834(n250 ,n14[1] ,n14[0]);
    not g835(n249 ,n14[1]);
    not g836(n248 ,n14[0]);
    not g837(n848 ,n1);
    nor g838(n849 ,n848 ,n847);
    or g839(n847 ,n844 ,n846);
    nor g840(n846 ,n845 ,n843);
    or g841(n845 ,n841 ,n842);
    nor g842(n844 ,n2[13] ,n2[12]);
    nor g843(n843 ,n2[11] ,n2[10]);
    not g844(n842 ,n2[12]);
    not g845(n841 ,n2[13]);
    nor g846(n11[11] ,n839 ,n840);
    nor g847(n840 ,n806 ,n838);
    nor g848(n839 ,n3[11] ,n837);
    nor g849(n11[10] ,n836 ,n837);
    not g850(n838 ,n837);
    nor g851(n837 ,n799 ,n835);
    nor g852(n836 ,n3[10] ,n834);
    nor g853(n11[9] ,n833 ,n834);
    not g854(n835 ,n834);
    nor g855(n834 ,n800 ,n832);
    nor g856(n833 ,n3[9] ,n831);
    nor g857(n11[8] ,n830 ,n831);
    not g858(n832 ,n831);
    nor g859(n831 ,n804 ,n829);
    nor g860(n830 ,n3[8] ,n828);
    nor g861(n11[7] ,n827 ,n828);
    not g862(n829 ,n828);
    nor g863(n828 ,n798 ,n826);
    nor g864(n827 ,n3[7] ,n825);
    nor g865(n11[6] ,n824 ,n825);
    not g866(n826 ,n825);
    nor g867(n825 ,n803 ,n823);
    nor g868(n824 ,n3[6] ,n822);
    nor g869(n11[5] ,n821 ,n822);
    not g870(n823 ,n822);
    nor g871(n822 ,n801 ,n820);
    nor g872(n821 ,n3[5] ,n819);
    nor g873(n11[4] ,n818 ,n819);
    not g874(n820 ,n819);
    nor g875(n819 ,n802 ,n817);
    nor g876(n818 ,n3[4] ,n816);
    nor g877(n11[3] ,n815 ,n816);
    not g878(n817 ,n816);
    nor g879(n816 ,n807 ,n814);
    nor g880(n815 ,n3[3] ,n813);
    nor g881(n11[2] ,n812 ,n813);
    not g882(n814 ,n813);
    nor g883(n813 ,n808 ,n811);
    nor g884(n812 ,n3[2] ,n810);
    nor g885(n11[1] ,n810 ,n809);
    not g886(n811 ,n810);
    nor g887(n810 ,n797 ,n805);
    nor g888(n809 ,n3[1] ,n849);
    not g889(n808 ,n3[2]);
    not g890(n807 ,n3[3]);
    not g891(n806 ,n3[11]);
    not g892(n805 ,n849);
    not g893(n804 ,n3[8]);
    not g894(n803 ,n3[6]);
    not g895(n802 ,n3[4]);
    not g896(n801 ,n3[5]);
    not g897(n800 ,n3[9]);
    not g898(n799 ,n3[10]);
    not g899(n798 ,n3[7]);
    not g900(n797 ,n3[1]);
endmodule
